module dadda_mult(
    output wire [63:0] Product,
    input wire [31:0] A,
    input wire [31:0] B
);

// Stage 0 partial products
wire[0:0] p_0_0; wire[1:0] p_0_1; wire[2:0] p_0_2; wire[3:0] p_0_3; wire[4:0] p_0_4; wire[5:0] p_0_5; wire[6:0] p_0_6; wire[7:0] p_0_7; wire[8:0] p_0_8; wire[9:0] p_0_9; wire[10:0] p_0_10; wire[11:0] p_0_11; wire[12:0] p_0_12; wire[13:0] p_0_13; wire[14:0] p_0_14; wire[15:0] p_0_15; wire[16:0] p_0_16; wire[17:0] p_0_17; wire[18:0] p_0_18; wire[19:0] p_0_19; wire[20:0] p_0_20; wire[21:0] p_0_21; wire[22:0] p_0_22; wire[23:0] p_0_23; wire[24:0] p_0_24; wire[25:0] p_0_25; wire[26:0] p_0_26; wire[27:0] p_0_27; wire[28:0] p_0_28; wire[29:0] p_0_29; wire[30:0] p_0_30; wire[31:0] p_0_31; wire[30:0] p_0_32; wire[29:0] p_0_33; wire[28:0] p_0_34; wire[27:0] p_0_35; wire[26:0] p_0_36; wire[25:0] p_0_37; wire[24:0] p_0_38; wire[23:0] p_0_39; wire[22:0] p_0_40; wire[21:0] p_0_41; wire[20:0] p_0_42; wire[19:0] p_0_43; wire[18:0] p_0_44; wire[17:0] p_0_45; wire[16:0] p_0_46; wire[15:0] p_0_47; wire[14:0] p_0_48; wire[13:0] p_0_49; wire[12:0] p_0_50; wire[11:0] p_0_51; wire[10:0] p_0_52; wire[9:0] p_0_53; wire[8:0] p_0_54; wire[7:0] p_0_55; wire[6:0] p_0_56; wire[5:0] p_0_57; wire[4:0] p_0_58; wire[3:0] p_0_59; wire[2:0] p_0_60; wire[1:0] p_0_61; wire[0:0] p_0_62; 
// Stage 1 partial products
wire[0:0] p_1_0; wire[1:0] p_1_1; wire[2:0] p_1_2; wire[3:0] p_1_3; wire[4:0] p_1_4; wire[5:0] p_1_5; wire[6:0] p_1_6; wire[7:0] p_1_7; wire[8:0] p_1_8; wire[9:0] p_1_9; wire[10:0] p_1_10; wire[11:0] p_1_11; wire[12:0] p_1_12; wire[13:0] p_1_13; wire[14:0] p_1_14; wire[15:0] p_1_15; wire[16:0] p_1_16; wire[17:0] p_1_17; wire[18:0] p_1_18; wire[19:0] p_1_19; wire[20:0] p_1_20; wire[21:0] p_1_21; wire[22:0] p_1_22; wire[23:0] p_1_23; wire[24:0] p_1_24; wire[25:0] p_1_25; wire[26:0] p_1_26; wire[27:0] p_1_27; wire[27:0] p_1_28; wire[27:0] p_1_29; wire[27:0] p_1_30; wire[27:0] p_1_31; wire[27:0] p_1_32; wire[27:0] p_1_33; wire[27:0] p_1_34; wire[27:0] p_1_35; wire[27:0] p_1_36; wire[25:0] p_1_37; wire[24:0] p_1_38; wire[23:0] p_1_39; wire[22:0] p_1_40; wire[21:0] p_1_41; wire[20:0] p_1_42; wire[19:0] p_1_43; wire[18:0] p_1_44; wire[17:0] p_1_45; wire[16:0] p_1_46; wire[15:0] p_1_47; wire[14:0] p_1_48; wire[13:0] p_1_49; wire[12:0] p_1_50; wire[11:0] p_1_51; wire[10:0] p_1_52; wire[9:0] p_1_53; wire[8:0] p_1_54; wire[7:0] p_1_55; wire[6:0] p_1_56; wire[5:0] p_1_57; wire[4:0] p_1_58; wire[3:0] p_1_59; wire[2:0] p_1_60; wire[1:0] p_1_61; wire[0:0] p_1_62; 
// Stage 2 partial products
wire[0:0] p_2_0; wire[1:0] p_2_1; wire[2:0] p_2_2; wire[3:0] p_2_3; wire[4:0] p_2_4; wire[5:0] p_2_5; wire[6:0] p_2_6; wire[7:0] p_2_7; wire[8:0] p_2_8; wire[9:0] p_2_9; wire[10:0] p_2_10; wire[11:0] p_2_11; wire[12:0] p_2_12; wire[13:0] p_2_13; wire[14:0] p_2_14; wire[15:0] p_2_15; wire[16:0] p_2_16; wire[17:0] p_2_17; wire[18:0] p_2_18; wire[18:0] p_2_19; wire[18:0] p_2_20; wire[18:0] p_2_21; wire[18:0] p_2_22; wire[18:0] p_2_23; wire[18:0] p_2_24; wire[18:0] p_2_25; wire[18:0] p_2_26; wire[18:0] p_2_27; wire[18:0] p_2_28; wire[18:0] p_2_29; wire[18:0] p_2_30; wire[18:0] p_2_31; wire[18:0] p_2_32; wire[18:0] p_2_33; wire[18:0] p_2_34; wire[18:0] p_2_35; wire[18:0] p_2_36; wire[18:0] p_2_37; wire[18:0] p_2_38; wire[18:0] p_2_39; wire[18:0] p_2_40; wire[18:0] p_2_41; wire[18:0] p_2_42; wire[18:0] p_2_43; wire[18:0] p_2_44; wire[18:0] p_2_45; wire[16:0] p_2_46; wire[15:0] p_2_47; wire[14:0] p_2_48; wire[13:0] p_2_49; wire[12:0] p_2_50; wire[11:0] p_2_51; wire[10:0] p_2_52; wire[9:0] p_2_53; wire[8:0] p_2_54; wire[7:0] p_2_55; wire[6:0] p_2_56; wire[5:0] p_2_57; wire[4:0] p_2_58; wire[3:0] p_2_59; wire[2:0] p_2_60; wire[1:0] p_2_61; wire[0:0] p_2_62; 
// Stage 3 partial products
wire[0:0] p_3_0; wire[1:0] p_3_1; wire[2:0] p_3_2; wire[3:0] p_3_3; wire[4:0] p_3_4; wire[5:0] p_3_5; wire[6:0] p_3_6; wire[7:0] p_3_7; wire[8:0] p_3_8; wire[9:0] p_3_9; wire[10:0] p_3_10; wire[11:0] p_3_11; wire[12:0] p_3_12; wire[12:0] p_3_13; wire[12:0] p_3_14; wire[12:0] p_3_15; wire[12:0] p_3_16; wire[12:0] p_3_17; wire[12:0] p_3_18; wire[12:0] p_3_19; wire[12:0] p_3_20; wire[12:0] p_3_21; wire[12:0] p_3_22; wire[12:0] p_3_23; wire[12:0] p_3_24; wire[12:0] p_3_25; wire[12:0] p_3_26; wire[12:0] p_3_27; wire[12:0] p_3_28; wire[12:0] p_3_29; wire[12:0] p_3_30; wire[12:0] p_3_31; wire[12:0] p_3_32; wire[12:0] p_3_33; wire[12:0] p_3_34; wire[12:0] p_3_35; wire[12:0] p_3_36; wire[12:0] p_3_37; wire[12:0] p_3_38; wire[12:0] p_3_39; wire[12:0] p_3_40; wire[12:0] p_3_41; wire[12:0] p_3_42; wire[12:0] p_3_43; wire[12:0] p_3_44; wire[12:0] p_3_45; wire[12:0] p_3_46; wire[12:0] p_3_47; wire[12:0] p_3_48; wire[12:0] p_3_49; wire[12:0] p_3_50; wire[12:0] p_3_51; wire[10:0] p_3_52; wire[9:0] p_3_53; wire[8:0] p_3_54; wire[7:0] p_3_55; wire[6:0] p_3_56; wire[5:0] p_3_57; wire[4:0] p_3_58; wire[3:0] p_3_59; wire[2:0] p_3_60; wire[1:0] p_3_61; wire[0:0] p_3_62; 
// Stage 4 partial products
wire[0:0] p_4_0; wire[1:0] p_4_1; wire[2:0] p_4_2; wire[3:0] p_4_3; wire[4:0] p_4_4; wire[5:0] p_4_5; wire[6:0] p_4_6; wire[7:0] p_4_7; wire[8:0] p_4_8; wire[8:0] p_4_9; wire[8:0] p_4_10; wire[8:0] p_4_11; wire[8:0] p_4_12; wire[8:0] p_4_13; wire[8:0] p_4_14; wire[8:0] p_4_15; wire[8:0] p_4_16; wire[8:0] p_4_17; wire[8:0] p_4_18; wire[8:0] p_4_19; wire[8:0] p_4_20; wire[8:0] p_4_21; wire[8:0] p_4_22; wire[8:0] p_4_23; wire[8:0] p_4_24; wire[8:0] p_4_25; wire[8:0] p_4_26; wire[8:0] p_4_27; wire[8:0] p_4_28; wire[8:0] p_4_29; wire[8:0] p_4_30; wire[8:0] p_4_31; wire[8:0] p_4_32; wire[8:0] p_4_33; wire[8:0] p_4_34; wire[8:0] p_4_35; wire[8:0] p_4_36; wire[8:0] p_4_37; wire[8:0] p_4_38; wire[8:0] p_4_39; wire[8:0] p_4_40; wire[8:0] p_4_41; wire[8:0] p_4_42; wire[8:0] p_4_43; wire[8:0] p_4_44; wire[8:0] p_4_45; wire[8:0] p_4_46; wire[8:0] p_4_47; wire[8:0] p_4_48; wire[8:0] p_4_49; wire[8:0] p_4_50; wire[8:0] p_4_51; wire[8:0] p_4_52; wire[8:0] p_4_53; wire[8:0] p_4_54; wire[8:0] p_4_55; wire[6:0] p_4_56; wire[5:0] p_4_57; wire[4:0] p_4_58; wire[3:0] p_4_59; wire[2:0] p_4_60; wire[1:0] p_4_61; wire[0:0] p_4_62; 
// Stage 5 partial products
wire[0:0] p_5_0; wire[1:0] p_5_1; wire[2:0] p_5_2; wire[3:0] p_5_3; wire[4:0] p_5_4; wire[5:0] p_5_5; wire[5:0] p_5_6; wire[5:0] p_5_7; wire[5:0] p_5_8; wire[5:0] p_5_9; wire[5:0] p_5_10; wire[5:0] p_5_11; wire[5:0] p_5_12; wire[5:0] p_5_13; wire[5:0] p_5_14; wire[5:0] p_5_15; wire[5:0] p_5_16; wire[5:0] p_5_17; wire[5:0] p_5_18; wire[5:0] p_5_19; wire[5:0] p_5_20; wire[5:0] p_5_21; wire[5:0] p_5_22; wire[5:0] p_5_23; wire[5:0] p_5_24; wire[5:0] p_5_25; wire[5:0] p_5_26; wire[5:0] p_5_27; wire[5:0] p_5_28; wire[5:0] p_5_29; wire[5:0] p_5_30; wire[5:0] p_5_31; wire[5:0] p_5_32; wire[5:0] p_5_33; wire[5:0] p_5_34; wire[5:0] p_5_35; wire[5:0] p_5_36; wire[5:0] p_5_37; wire[5:0] p_5_38; wire[5:0] p_5_39; wire[5:0] p_5_40; wire[5:0] p_5_41; wire[5:0] p_5_42; wire[5:0] p_5_43; wire[5:0] p_5_44; wire[5:0] p_5_45; wire[5:0] p_5_46; wire[5:0] p_5_47; wire[5:0] p_5_48; wire[5:0] p_5_49; wire[5:0] p_5_50; wire[5:0] p_5_51; wire[5:0] p_5_52; wire[5:0] p_5_53; wire[5:0] p_5_54; wire[5:0] p_5_55; wire[5:0] p_5_56; wire[5:0] p_5_57; wire[5:0] p_5_58; wire[3:0] p_5_59; wire[2:0] p_5_60; wire[1:0] p_5_61; wire[0:0] p_5_62; 
// Stage 6 partial products
wire[0:0] p_6_0; wire[1:0] p_6_1; wire[2:0] p_6_2; wire[3:0] p_6_3; wire[3:0] p_6_4; wire[3:0] p_6_5; wire[3:0] p_6_6; wire[3:0] p_6_7; wire[3:0] p_6_8; wire[3:0] p_6_9; wire[3:0] p_6_10; wire[3:0] p_6_11; wire[3:0] p_6_12; wire[3:0] p_6_13; wire[3:0] p_6_14; wire[3:0] p_6_15; wire[3:0] p_6_16; wire[3:0] p_6_17; wire[3:0] p_6_18; wire[3:0] p_6_19; wire[3:0] p_6_20; wire[3:0] p_6_21; wire[3:0] p_6_22; wire[3:0] p_6_23; wire[3:0] p_6_24; wire[3:0] p_6_25; wire[3:0] p_6_26; wire[3:0] p_6_27; wire[3:0] p_6_28; wire[3:0] p_6_29; wire[3:0] p_6_30; wire[3:0] p_6_31; wire[3:0] p_6_32; wire[3:0] p_6_33; wire[3:0] p_6_34; wire[3:0] p_6_35; wire[3:0] p_6_36; wire[3:0] p_6_37; wire[3:0] p_6_38; wire[3:0] p_6_39; wire[3:0] p_6_40; wire[3:0] p_6_41; wire[3:0] p_6_42; wire[3:0] p_6_43; wire[3:0] p_6_44; wire[3:0] p_6_45; wire[3:0] p_6_46; wire[3:0] p_6_47; wire[3:0] p_6_48; wire[3:0] p_6_49; wire[3:0] p_6_50; wire[3:0] p_6_51; wire[3:0] p_6_52; wire[3:0] p_6_53; wire[3:0] p_6_54; wire[3:0] p_6_55; wire[3:0] p_6_56; wire[3:0] p_6_57; wire[3:0] p_6_58; wire[3:0] p_6_59; wire[3:0] p_6_60; wire[1:0] p_6_61; wire[0:0] p_6_62; 
// Stage 7 partial products
wire[0:0] p_7_0; wire[1:0] p_7_1; wire[2:0] p_7_2; wire[2:0] p_7_3; wire[2:0] p_7_4; wire[2:0] p_7_5; wire[2:0] p_7_6; wire[2:0] p_7_7; wire[2:0] p_7_8; wire[2:0] p_7_9; wire[2:0] p_7_10; wire[2:0] p_7_11; wire[2:0] p_7_12; wire[2:0] p_7_13; wire[2:0] p_7_14; wire[2:0] p_7_15; wire[2:0] p_7_16; wire[2:0] p_7_17; wire[2:0] p_7_18; wire[2:0] p_7_19; wire[2:0] p_7_20; wire[2:0] p_7_21; wire[2:0] p_7_22; wire[2:0] p_7_23; wire[2:0] p_7_24; wire[2:0] p_7_25; wire[2:0] p_7_26; wire[2:0] p_7_27; wire[2:0] p_7_28; wire[2:0] p_7_29; wire[2:0] p_7_30; wire[2:0] p_7_31; wire[2:0] p_7_32; wire[2:0] p_7_33; wire[2:0] p_7_34; wire[2:0] p_7_35; wire[2:0] p_7_36; wire[2:0] p_7_37; wire[2:0] p_7_38; wire[2:0] p_7_39; wire[2:0] p_7_40; wire[2:0] p_7_41; wire[2:0] p_7_42; wire[2:0] p_7_43; wire[2:0] p_7_44; wire[2:0] p_7_45; wire[2:0] p_7_46; wire[2:0] p_7_47; wire[2:0] p_7_48; wire[2:0] p_7_49; wire[2:0] p_7_50; wire[2:0] p_7_51; wire[2:0] p_7_52; wire[2:0] p_7_53; wire[2:0] p_7_54; wire[2:0] p_7_55; wire[2:0] p_7_56; wire[2:0] p_7_57; wire[2:0] p_7_58; wire[2:0] p_7_59; wire[2:0] p_7_60; wire[2:0] p_7_61; wire[0:0] p_7_62; 
// Stage 8 partial products
wire[0:0] p_8_0; wire[1:0] p_8_1; wire[1:0] p_8_2; wire[1:0] p_8_3; wire[1:0] p_8_4; wire[1:0] p_8_5; wire[1:0] p_8_6; wire[1:0] p_8_7; wire[1:0] p_8_8; wire[1:0] p_8_9; wire[1:0] p_8_10; wire[1:0] p_8_11; wire[1:0] p_8_12; wire[1:0] p_8_13; wire[1:0] p_8_14; wire[1:0] p_8_15; wire[1:0] p_8_16; wire[1:0] p_8_17; wire[1:0] p_8_18; wire[1:0] p_8_19; wire[1:0] p_8_20; wire[1:0] p_8_21; wire[1:0] p_8_22; wire[1:0] p_8_23; wire[1:0] p_8_24; wire[1:0] p_8_25; wire[1:0] p_8_26; wire[1:0] p_8_27; wire[1:0] p_8_28; wire[1:0] p_8_29; wire[1:0] p_8_30; wire[1:0] p_8_31; wire[1:0] p_8_32; wire[1:0] p_8_33; wire[1:0] p_8_34; wire[1:0] p_8_35; wire[1:0] p_8_36; wire[1:0] p_8_37; wire[1:0] p_8_38; wire[1:0] p_8_39; wire[1:0] p_8_40; wire[1:0] p_8_41; wire[1:0] p_8_42; wire[1:0] p_8_43; wire[1:0] p_8_44; wire[1:0] p_8_45; wire[1:0] p_8_46; wire[1:0] p_8_47; wire[1:0] p_8_48; wire[1:0] p_8_49; wire[1:0] p_8_50; wire[1:0] p_8_51; wire[1:0] p_8_52; wire[1:0] p_8_53; wire[1:0] p_8_54; wire[1:0] p_8_55; wire[1:0] p_8_56; wire[1:0] p_8_57; wire[1:0] p_8_58; wire[1:0] p_8_59; wire[1:0] p_8_60; wire[1:0] p_8_61; wire[1:0] p_8_62; 

// AND gate array
assign p_0_0 = {A[0]&B[0]};
assign p_0_1 = {A[1]&B[0], A[0]&B[1]};
assign p_0_2 = {A[2]&B[0], A[1]&B[1], A[0]&B[2]};
assign p_0_3 = {A[3]&B[0], A[2]&B[1], A[1]&B[2], A[0]&B[3]};
assign p_0_4 = {A[4]&B[0], A[3]&B[1], A[2]&B[2], A[1]&B[3], A[0]&B[4]};
assign p_0_5 = {A[5]&B[0], A[4]&B[1], A[3]&B[2], A[2]&B[3], A[1]&B[4], A[0]&B[5]};
assign p_0_6 = {A[6]&B[0], A[5]&B[1], A[4]&B[2], A[3]&B[3], A[2]&B[4], A[1]&B[5], A[0]&B[6]};
assign p_0_7 = {A[7]&B[0], A[6]&B[1], A[5]&B[2], A[4]&B[3], A[3]&B[4], A[2]&B[5], A[1]&B[6], A[0]&B[7]};
assign p_0_8 = {A[8]&B[0], A[7]&B[1], A[6]&B[2], A[5]&B[3], A[4]&B[4], A[3]&B[5], A[2]&B[6], A[1]&B[7], A[0]&B[8]};
assign p_0_9 = {A[9]&B[0], A[8]&B[1], A[7]&B[2], A[6]&B[3], A[5]&B[4], A[4]&B[5], A[3]&B[6], A[2]&B[7], A[1]&B[8], A[0]&B[9]};
assign p_0_10 = {A[10]&B[0], A[9]&B[1], A[8]&B[2], A[7]&B[3], A[6]&B[4], A[5]&B[5], A[4]&B[6], A[3]&B[7], A[2]&B[8], A[1]&B[9], A[0]&B[10]};
assign p_0_11 = {A[11]&B[0], A[10]&B[1], A[9]&B[2], A[8]&B[3], A[7]&B[4], A[6]&B[5], A[5]&B[6], A[4]&B[7], A[3]&B[8], A[2]&B[9], A[1]&B[10], A[0]&B[11]};
assign p_0_12 = {A[12]&B[0], A[11]&B[1], A[10]&B[2], A[9]&B[3], A[8]&B[4], A[7]&B[5], A[6]&B[6], A[5]&B[7], A[4]&B[8], A[3]&B[9], A[2]&B[10], A[1]&B[11], A[0]&B[12]};
assign p_0_13 = {A[13]&B[0], A[12]&B[1], A[11]&B[2], A[10]&B[3], A[9]&B[4], A[8]&B[5], A[7]&B[6], A[6]&B[7], A[5]&B[8], A[4]&B[9], A[3]&B[10], A[2]&B[11], A[1]&B[12], A[0]&B[13]};
assign p_0_14 = {A[14]&B[0], A[13]&B[1], A[12]&B[2], A[11]&B[3], A[10]&B[4], A[9]&B[5], A[8]&B[6], A[7]&B[7], A[6]&B[8], A[5]&B[9], A[4]&B[10], A[3]&B[11], A[2]&B[12], A[1]&B[13], A[0]&B[14]};
assign p_0_15 = {A[15]&B[0], A[14]&B[1], A[13]&B[2], A[12]&B[3], A[11]&B[4], A[10]&B[5], A[9]&B[6], A[8]&B[7], A[7]&B[8], A[6]&B[9], A[5]&B[10], A[4]&B[11], A[3]&B[12], A[2]&B[13], A[1]&B[14], A[0]&B[15]};
assign p_0_16 = {A[16]&B[0], A[15]&B[1], A[14]&B[2], A[13]&B[3], A[12]&B[4], A[11]&B[5], A[10]&B[6], A[9]&B[7], A[8]&B[8], A[7]&B[9], A[6]&B[10], A[5]&B[11], A[4]&B[12], A[3]&B[13], A[2]&B[14], A[1]&B[15], A[0]&B[16]};
assign p_0_17 = {A[17]&B[0], A[16]&B[1], A[15]&B[2], A[14]&B[3], A[13]&B[4], A[12]&B[5], A[11]&B[6], A[10]&B[7], A[9]&B[8], A[8]&B[9], A[7]&B[10], A[6]&B[11], A[5]&B[12], A[4]&B[13], A[3]&B[14], A[2]&B[15], A[1]&B[16], A[0]&B[17]};
assign p_0_18 = {A[18]&B[0], A[17]&B[1], A[16]&B[2], A[15]&B[3], A[14]&B[4], A[13]&B[5], A[12]&B[6], A[11]&B[7], A[10]&B[8], A[9]&B[9], A[8]&B[10], A[7]&B[11], A[6]&B[12], A[5]&B[13], A[4]&B[14], A[3]&B[15], A[2]&B[16], A[1]&B[17], A[0]&B[18]};
assign p_0_19 = {A[19]&B[0], A[18]&B[1], A[17]&B[2], A[16]&B[3], A[15]&B[4], A[14]&B[5], A[13]&B[6], A[12]&B[7], A[11]&B[8], A[10]&B[9], A[9]&B[10], A[8]&B[11], A[7]&B[12], A[6]&B[13], A[5]&B[14], A[4]&B[15], A[3]&B[16], A[2]&B[17], A[1]&B[18], A[0]&B[19]};
assign p_0_20 = {A[20]&B[0], A[19]&B[1], A[18]&B[2], A[17]&B[3], A[16]&B[4], A[15]&B[5], A[14]&B[6], A[13]&B[7], A[12]&B[8], A[11]&B[9], A[10]&B[10], A[9]&B[11], A[8]&B[12], A[7]&B[13], A[6]&B[14], A[5]&B[15], A[4]&B[16], A[3]&B[17], A[2]&B[18], A[1]&B[19], A[0]&B[20]};
assign p_0_21 = {A[21]&B[0], A[20]&B[1], A[19]&B[2], A[18]&B[3], A[17]&B[4], A[16]&B[5], A[15]&B[6], A[14]&B[7], A[13]&B[8], A[12]&B[9], A[11]&B[10], A[10]&B[11], A[9]&B[12], A[8]&B[13], A[7]&B[14], A[6]&B[15], A[5]&B[16], A[4]&B[17], A[3]&B[18], A[2]&B[19], A[1]&B[20], A[0]&B[21]};
assign p_0_22 = {A[22]&B[0], A[21]&B[1], A[20]&B[2], A[19]&B[3], A[18]&B[4], A[17]&B[5], A[16]&B[6], A[15]&B[7], A[14]&B[8], A[13]&B[9], A[12]&B[10], A[11]&B[11], A[10]&B[12], A[9]&B[13], A[8]&B[14], A[7]&B[15], A[6]&B[16], A[5]&B[17], A[4]&B[18], A[3]&B[19], A[2]&B[20], A[1]&B[21], A[0]&B[22]};
assign p_0_23 = {A[23]&B[0], A[22]&B[1], A[21]&B[2], A[20]&B[3], A[19]&B[4], A[18]&B[5], A[17]&B[6], A[16]&B[7], A[15]&B[8], A[14]&B[9], A[13]&B[10], A[12]&B[11], A[11]&B[12], A[10]&B[13], A[9]&B[14], A[8]&B[15], A[7]&B[16], A[6]&B[17], A[5]&B[18], A[4]&B[19], A[3]&B[20], A[2]&B[21], A[1]&B[22], A[0]&B[23]};
assign p_0_24 = {A[24]&B[0], A[23]&B[1], A[22]&B[2], A[21]&B[3], A[20]&B[4], A[19]&B[5], A[18]&B[6], A[17]&B[7], A[16]&B[8], A[15]&B[9], A[14]&B[10], A[13]&B[11], A[12]&B[12], A[11]&B[13], A[10]&B[14], A[9]&B[15], A[8]&B[16], A[7]&B[17], A[6]&B[18], A[5]&B[19], A[4]&B[20], A[3]&B[21], A[2]&B[22], A[1]&B[23], A[0]&B[24]};
assign p_0_25 = {A[25]&B[0], A[24]&B[1], A[23]&B[2], A[22]&B[3], A[21]&B[4], A[20]&B[5], A[19]&B[6], A[18]&B[7], A[17]&B[8], A[16]&B[9], A[15]&B[10], A[14]&B[11], A[13]&B[12], A[12]&B[13], A[11]&B[14], A[10]&B[15], A[9]&B[16], A[8]&B[17], A[7]&B[18], A[6]&B[19], A[5]&B[20], A[4]&B[21], A[3]&B[22], A[2]&B[23], A[1]&B[24], A[0]&B[25]};
assign p_0_26 = {A[26]&B[0], A[25]&B[1], A[24]&B[2], A[23]&B[3], A[22]&B[4], A[21]&B[5], A[20]&B[6], A[19]&B[7], A[18]&B[8], A[17]&B[9], A[16]&B[10], A[15]&B[11], A[14]&B[12], A[13]&B[13], A[12]&B[14], A[11]&B[15], A[10]&B[16], A[9]&B[17], A[8]&B[18], A[7]&B[19], A[6]&B[20], A[5]&B[21], A[4]&B[22], A[3]&B[23], A[2]&B[24], A[1]&B[25], A[0]&B[26]};
assign p_0_27 = {A[27]&B[0], A[26]&B[1], A[25]&B[2], A[24]&B[3], A[23]&B[4], A[22]&B[5], A[21]&B[6], A[20]&B[7], A[19]&B[8], A[18]&B[9], A[17]&B[10], A[16]&B[11], A[15]&B[12], A[14]&B[13], A[13]&B[14], A[12]&B[15], A[11]&B[16], A[10]&B[17], A[9]&B[18], A[8]&B[19], A[7]&B[20], A[6]&B[21], A[5]&B[22], A[4]&B[23], A[3]&B[24], A[2]&B[25], A[1]&B[26], A[0]&B[27]};
assign p_0_28 = {A[28]&B[0], A[27]&B[1], A[26]&B[2], A[25]&B[3], A[24]&B[4], A[23]&B[5], A[22]&B[6], A[21]&B[7], A[20]&B[8], A[19]&B[9], A[18]&B[10], A[17]&B[11], A[16]&B[12], A[15]&B[13], A[14]&B[14], A[13]&B[15], A[12]&B[16], A[11]&B[17], A[10]&B[18], A[9]&B[19], A[8]&B[20], A[7]&B[21], A[6]&B[22], A[5]&B[23], A[4]&B[24], A[3]&B[25], A[2]&B[26], A[1]&B[27], A[0]&B[28]};
assign p_0_29 = {A[29]&B[0], A[28]&B[1], A[27]&B[2], A[26]&B[3], A[25]&B[4], A[24]&B[5], A[23]&B[6], A[22]&B[7], A[21]&B[8], A[20]&B[9], A[19]&B[10], A[18]&B[11], A[17]&B[12], A[16]&B[13], A[15]&B[14], A[14]&B[15], A[13]&B[16], A[12]&B[17], A[11]&B[18], A[10]&B[19], A[9]&B[20], A[8]&B[21], A[7]&B[22], A[6]&B[23], A[5]&B[24], A[4]&B[25], A[3]&B[26], A[2]&B[27], A[1]&B[28], A[0]&B[29]};
assign p_0_30 = {A[30]&B[0], A[29]&B[1], A[28]&B[2], A[27]&B[3], A[26]&B[4], A[25]&B[5], A[24]&B[6], A[23]&B[7], A[22]&B[8], A[21]&B[9], A[20]&B[10], A[19]&B[11], A[18]&B[12], A[17]&B[13], A[16]&B[14], A[15]&B[15], A[14]&B[16], A[13]&B[17], A[12]&B[18], A[11]&B[19], A[10]&B[20], A[9]&B[21], A[8]&B[22], A[7]&B[23], A[6]&B[24], A[5]&B[25], A[4]&B[26], A[3]&B[27], A[2]&B[28], A[1]&B[29], A[0]&B[30]};
assign p_0_31 = {A[31]&B[0], A[30]&B[1], A[29]&B[2], A[28]&B[3], A[27]&B[4], A[26]&B[5], A[25]&B[6], A[24]&B[7], A[23]&B[8], A[22]&B[9], A[21]&B[10], A[20]&B[11], A[19]&B[12], A[18]&B[13], A[17]&B[14], A[16]&B[15], A[15]&B[16], A[14]&B[17], A[13]&B[18], A[12]&B[19], A[11]&B[20], A[10]&B[21], A[9]&B[22], A[8]&B[23], A[7]&B[24], A[6]&B[25], A[5]&B[26], A[4]&B[27], A[3]&B[28], A[2]&B[29], A[1]&B[30], A[0]&B[31]};
assign p_0_32 = {A[31]&B[1], A[30]&B[2], A[29]&B[3], A[28]&B[4], A[27]&B[5], A[26]&B[6], A[25]&B[7], A[24]&B[8], A[23]&B[9], A[22]&B[10], A[21]&B[11], A[20]&B[12], A[19]&B[13], A[18]&B[14], A[17]&B[15], A[16]&B[16], A[15]&B[17], A[14]&B[18], A[13]&B[19], A[12]&B[20], A[11]&B[21], A[10]&B[22], A[9]&B[23], A[8]&B[24], A[7]&B[25], A[6]&B[26], A[5]&B[27], A[4]&B[28], A[3]&B[29], A[2]&B[30], A[1]&B[31]};
assign p_0_33 = {A[31]&B[2], A[30]&B[3], A[29]&B[4], A[28]&B[5], A[27]&B[6], A[26]&B[7], A[25]&B[8], A[24]&B[9], A[23]&B[10], A[22]&B[11], A[21]&B[12], A[20]&B[13], A[19]&B[14], A[18]&B[15], A[17]&B[16], A[16]&B[17], A[15]&B[18], A[14]&B[19], A[13]&B[20], A[12]&B[21], A[11]&B[22], A[10]&B[23], A[9]&B[24], A[8]&B[25], A[7]&B[26], A[6]&B[27], A[5]&B[28], A[4]&B[29], A[3]&B[30], A[2]&B[31]};
assign p_0_34 = {A[31]&B[3], A[30]&B[4], A[29]&B[5], A[28]&B[6], A[27]&B[7], A[26]&B[8], A[25]&B[9], A[24]&B[10], A[23]&B[11], A[22]&B[12], A[21]&B[13], A[20]&B[14], A[19]&B[15], A[18]&B[16], A[17]&B[17], A[16]&B[18], A[15]&B[19], A[14]&B[20], A[13]&B[21], A[12]&B[22], A[11]&B[23], A[10]&B[24], A[9]&B[25], A[8]&B[26], A[7]&B[27], A[6]&B[28], A[5]&B[29], A[4]&B[30], A[3]&B[31]};
assign p_0_35 = {A[31]&B[4], A[30]&B[5], A[29]&B[6], A[28]&B[7], A[27]&B[8], A[26]&B[9], A[25]&B[10], A[24]&B[11], A[23]&B[12], A[22]&B[13], A[21]&B[14], A[20]&B[15], A[19]&B[16], A[18]&B[17], A[17]&B[18], A[16]&B[19], A[15]&B[20], A[14]&B[21], A[13]&B[22], A[12]&B[23], A[11]&B[24], A[10]&B[25], A[9]&B[26], A[8]&B[27], A[7]&B[28], A[6]&B[29], A[5]&B[30], A[4]&B[31]};
assign p_0_36 = {A[31]&B[5], A[30]&B[6], A[29]&B[7], A[28]&B[8], A[27]&B[9], A[26]&B[10], A[25]&B[11], A[24]&B[12], A[23]&B[13], A[22]&B[14], A[21]&B[15], A[20]&B[16], A[19]&B[17], A[18]&B[18], A[17]&B[19], A[16]&B[20], A[15]&B[21], A[14]&B[22], A[13]&B[23], A[12]&B[24], A[11]&B[25], A[10]&B[26], A[9]&B[27], A[8]&B[28], A[7]&B[29], A[6]&B[30], A[5]&B[31]};
assign p_0_37 = {A[31]&B[6], A[30]&B[7], A[29]&B[8], A[28]&B[9], A[27]&B[10], A[26]&B[11], A[25]&B[12], A[24]&B[13], A[23]&B[14], A[22]&B[15], A[21]&B[16], A[20]&B[17], A[19]&B[18], A[18]&B[19], A[17]&B[20], A[16]&B[21], A[15]&B[22], A[14]&B[23], A[13]&B[24], A[12]&B[25], A[11]&B[26], A[10]&B[27], A[9]&B[28], A[8]&B[29], A[7]&B[30], A[6]&B[31]};
assign p_0_38 = {A[31]&B[7], A[30]&B[8], A[29]&B[9], A[28]&B[10], A[27]&B[11], A[26]&B[12], A[25]&B[13], A[24]&B[14], A[23]&B[15], A[22]&B[16], A[21]&B[17], A[20]&B[18], A[19]&B[19], A[18]&B[20], A[17]&B[21], A[16]&B[22], A[15]&B[23], A[14]&B[24], A[13]&B[25], A[12]&B[26], A[11]&B[27], A[10]&B[28], A[9]&B[29], A[8]&B[30], A[7]&B[31]};
assign p_0_39 = {A[31]&B[8], A[30]&B[9], A[29]&B[10], A[28]&B[11], A[27]&B[12], A[26]&B[13], A[25]&B[14], A[24]&B[15], A[23]&B[16], A[22]&B[17], A[21]&B[18], A[20]&B[19], A[19]&B[20], A[18]&B[21], A[17]&B[22], A[16]&B[23], A[15]&B[24], A[14]&B[25], A[13]&B[26], A[12]&B[27], A[11]&B[28], A[10]&B[29], A[9]&B[30], A[8]&B[31]};
assign p_0_40 = {A[31]&B[9], A[30]&B[10], A[29]&B[11], A[28]&B[12], A[27]&B[13], A[26]&B[14], A[25]&B[15], A[24]&B[16], A[23]&B[17], A[22]&B[18], A[21]&B[19], A[20]&B[20], A[19]&B[21], A[18]&B[22], A[17]&B[23], A[16]&B[24], A[15]&B[25], A[14]&B[26], A[13]&B[27], A[12]&B[28], A[11]&B[29], A[10]&B[30], A[9]&B[31]};
assign p_0_41 = {A[31]&B[10], A[30]&B[11], A[29]&B[12], A[28]&B[13], A[27]&B[14], A[26]&B[15], A[25]&B[16], A[24]&B[17], A[23]&B[18], A[22]&B[19], A[21]&B[20], A[20]&B[21], A[19]&B[22], A[18]&B[23], A[17]&B[24], A[16]&B[25], A[15]&B[26], A[14]&B[27], A[13]&B[28], A[12]&B[29], A[11]&B[30], A[10]&B[31]};
assign p_0_42 = {A[31]&B[11], A[30]&B[12], A[29]&B[13], A[28]&B[14], A[27]&B[15], A[26]&B[16], A[25]&B[17], A[24]&B[18], A[23]&B[19], A[22]&B[20], A[21]&B[21], A[20]&B[22], A[19]&B[23], A[18]&B[24], A[17]&B[25], A[16]&B[26], A[15]&B[27], A[14]&B[28], A[13]&B[29], A[12]&B[30], A[11]&B[31]};
assign p_0_43 = {A[31]&B[12], A[30]&B[13], A[29]&B[14], A[28]&B[15], A[27]&B[16], A[26]&B[17], A[25]&B[18], A[24]&B[19], A[23]&B[20], A[22]&B[21], A[21]&B[22], A[20]&B[23], A[19]&B[24], A[18]&B[25], A[17]&B[26], A[16]&B[27], A[15]&B[28], A[14]&B[29], A[13]&B[30], A[12]&B[31]};
assign p_0_44 = {A[31]&B[13], A[30]&B[14], A[29]&B[15], A[28]&B[16], A[27]&B[17], A[26]&B[18], A[25]&B[19], A[24]&B[20], A[23]&B[21], A[22]&B[22], A[21]&B[23], A[20]&B[24], A[19]&B[25], A[18]&B[26], A[17]&B[27], A[16]&B[28], A[15]&B[29], A[14]&B[30], A[13]&B[31]};
assign p_0_45 = {A[31]&B[14], A[30]&B[15], A[29]&B[16], A[28]&B[17], A[27]&B[18], A[26]&B[19], A[25]&B[20], A[24]&B[21], A[23]&B[22], A[22]&B[23], A[21]&B[24], A[20]&B[25], A[19]&B[26], A[18]&B[27], A[17]&B[28], A[16]&B[29], A[15]&B[30], A[14]&B[31]};
assign p_0_46 = {A[31]&B[15], A[30]&B[16], A[29]&B[17], A[28]&B[18], A[27]&B[19], A[26]&B[20], A[25]&B[21], A[24]&B[22], A[23]&B[23], A[22]&B[24], A[21]&B[25], A[20]&B[26], A[19]&B[27], A[18]&B[28], A[17]&B[29], A[16]&B[30], A[15]&B[31]};
assign p_0_47 = {A[31]&B[16], A[30]&B[17], A[29]&B[18], A[28]&B[19], A[27]&B[20], A[26]&B[21], A[25]&B[22], A[24]&B[23], A[23]&B[24], A[22]&B[25], A[21]&B[26], A[20]&B[27], A[19]&B[28], A[18]&B[29], A[17]&B[30], A[16]&B[31]};
assign p_0_48 = {A[31]&B[17], A[30]&B[18], A[29]&B[19], A[28]&B[20], A[27]&B[21], A[26]&B[22], A[25]&B[23], A[24]&B[24], A[23]&B[25], A[22]&B[26], A[21]&B[27], A[20]&B[28], A[19]&B[29], A[18]&B[30], A[17]&B[31]};
assign p_0_49 = {A[31]&B[18], A[30]&B[19], A[29]&B[20], A[28]&B[21], A[27]&B[22], A[26]&B[23], A[25]&B[24], A[24]&B[25], A[23]&B[26], A[22]&B[27], A[21]&B[28], A[20]&B[29], A[19]&B[30], A[18]&B[31]};
assign p_0_50 = {A[31]&B[19], A[30]&B[20], A[29]&B[21], A[28]&B[22], A[27]&B[23], A[26]&B[24], A[25]&B[25], A[24]&B[26], A[23]&B[27], A[22]&B[28], A[21]&B[29], A[20]&B[30], A[19]&B[31]};
assign p_0_51 = {A[31]&B[20], A[30]&B[21], A[29]&B[22], A[28]&B[23], A[27]&B[24], A[26]&B[25], A[25]&B[26], A[24]&B[27], A[23]&B[28], A[22]&B[29], A[21]&B[30], A[20]&B[31]};
assign p_0_52 = {A[31]&B[21], A[30]&B[22], A[29]&B[23], A[28]&B[24], A[27]&B[25], A[26]&B[26], A[25]&B[27], A[24]&B[28], A[23]&B[29], A[22]&B[30], A[21]&B[31]};
assign p_0_53 = {A[31]&B[22], A[30]&B[23], A[29]&B[24], A[28]&B[25], A[27]&B[26], A[26]&B[27], A[25]&B[28], A[24]&B[29], A[23]&B[30], A[22]&B[31]};
assign p_0_54 = {A[31]&B[23], A[30]&B[24], A[29]&B[25], A[28]&B[26], A[27]&B[27], A[26]&B[28], A[25]&B[29], A[24]&B[30], A[23]&B[31]};
assign p_0_55 = {A[31]&B[24], A[30]&B[25], A[29]&B[26], A[28]&B[27], A[27]&B[28], A[26]&B[29], A[25]&B[30], A[24]&B[31]};
assign p_0_56 = {A[31]&B[25], A[30]&B[26], A[29]&B[27], A[28]&B[28], A[27]&B[29], A[26]&B[30], A[25]&B[31]};
assign p_0_57 = {A[31]&B[26], A[30]&B[27], A[29]&B[28], A[28]&B[29], A[27]&B[30], A[26]&B[31]};
assign p_0_58 = {A[31]&B[27], A[30]&B[28], A[29]&B[29], A[28]&B[30], A[27]&B[31]};
assign p_0_59 = {A[31]&B[28], A[30]&B[29], A[29]&B[30], A[28]&B[31]};
assign p_0_60 = {A[31]&B[29], A[30]&B[30], A[29]&B[31]};
assign p_0_61 = {A[31]&B[30], A[30]&B[31]};
assign p_0_62 = {A[31]&B[31]};

// Stage 1 non-added partial products
assign p_1_0[0:0] = p_0_0[0:0];
assign p_1_1[1:0] = p_0_1[1:0];
assign p_1_2[2:0] = p_0_2[2:0];
assign p_1_3[3:0] = p_0_3[3:0];
assign p_1_4[4:0] = p_0_4[4:0];
assign p_1_5[5:0] = p_0_5[5:0];
assign p_1_6[6:0] = p_0_6[6:0];
assign p_1_7[7:0] = p_0_7[7:0];
assign p_1_8[8:0] = p_0_8[8:0];
assign p_1_9[9:0] = p_0_9[9:0];
assign p_1_10[10:0] = p_0_10[10:0];
assign p_1_11[11:0] = p_0_11[11:0];
assign p_1_12[12:0] = p_0_12[12:0];
assign p_1_13[13:0] = p_0_13[13:0];
assign p_1_14[14:0] = p_0_14[14:0];
assign p_1_15[15:0] = p_0_15[15:0];
assign p_1_16[16:0] = p_0_16[16:0];
assign p_1_17[17:0] = p_0_17[17:0];
assign p_1_18[18:0] = p_0_18[18:0];
assign p_1_19[19:0] = p_0_19[19:0];
assign p_1_20[20:0] = p_0_20[20:0];
assign p_1_21[21:0] = p_0_21[21:0];
assign p_1_22[22:0] = p_0_22[22:0];
assign p_1_23[23:0] = p_0_23[23:0];
assign p_1_24[24:0] = p_0_24[24:0];
assign p_1_25[25:0] = p_0_25[25:0];
assign p_1_26[26:0] = p_0_26[26:0];
assign p_1_27[27:0] = p_0_27[27:0];
assign p_1_28[27:1] = p_0_28[26:0];
assign p_1_29[27:3] = p_0_29[24:0];
assign p_1_30[27:5] = p_0_30[22:0];
assign p_1_31[27:7] = p_0_31[20:0];
assign p_1_32[27:8] = p_0_32[19:0];
assign p_1_33[27:7] = p_0_33[20:0];
assign p_1_34[27:5] = p_0_34[22:0];
assign p_1_35[27:3] = p_0_35[24:0];
assign p_1_36[27:1] = p_0_36[26:0];
assign p_1_37[25:0] = p_0_37[25:0];
assign p_1_38[24:0] = p_0_38[24:0];
assign p_1_39[23:0] = p_0_39[23:0];
assign p_1_40[22:0] = p_0_40[22:0];
assign p_1_41[21:0] = p_0_41[21:0];
assign p_1_42[20:0] = p_0_42[20:0];
assign p_1_43[19:0] = p_0_43[19:0];
assign p_1_44[18:0] = p_0_44[18:0];
assign p_1_45[17:0] = p_0_45[17:0];
assign p_1_46[16:0] = p_0_46[16:0];
assign p_1_47[15:0] = p_0_47[15:0];
assign p_1_48[14:0] = p_0_48[14:0];
assign p_1_49[13:0] = p_0_49[13:0];
assign p_1_50[12:0] = p_0_50[12:0];
assign p_1_51[11:0] = p_0_51[11:0];
assign p_1_52[10:0] = p_0_52[10:0];
assign p_1_53[9:0] = p_0_53[9:0];
assign p_1_54[8:0] = p_0_54[8:0];
assign p_1_55[7:0] = p_0_55[7:0];
assign p_1_56[6:0] = p_0_56[6:0];
assign p_1_57[5:0] = p_0_57[5:0];
assign p_1_58[4:0] = p_0_58[4:0];
assign p_1_59[3:0] = p_0_59[3:0];
assign p_1_60[2:0] = p_0_60[2:0];
assign p_1_61[1:0] = p_0_61[1:0];
assign p_1_62[0:0] = p_0_62[0:0];
// Stage 1 adders
half_adder ha_1_28(.S(p_1_28[0]), .Cout(p_1_29[0]), .A(p_0_28[28]), .B(p_0_28[27]));
full_adder fa_1_29_0(.S(p_1_29[1]), .Cout(p_1_30[0]), .A(p_0_29[29]), .B(p_0_29[28]), .Cin(p_0_29[27]));
half_adder ha_1_29(.S(p_1_29[2]), .Cout(p_1_30[1]), .A(p_0_29[26]), .B(p_0_29[25]));
full_adder fa_1_30_0(.S(p_1_30[2]), .Cout(p_1_31[0]), .A(p_0_30[30]), .B(p_0_30[29]), .Cin(p_0_30[28]));
full_adder fa_1_30_1(.S(p_1_30[3]), .Cout(p_1_31[1]), .A(p_0_30[27]), .B(p_0_30[26]), .Cin(p_0_30[25]));
half_adder ha_1_30(.S(p_1_30[4]), .Cout(p_1_31[2]), .A(p_0_30[24]), .B(p_0_30[23]));
full_adder fa_1_31_0(.S(p_1_31[3]), .Cout(p_1_32[0]), .A(p_0_31[31]), .B(p_0_31[30]), .Cin(p_0_31[29]));
full_adder fa_1_31_1(.S(p_1_31[4]), .Cout(p_1_32[1]), .A(p_0_31[28]), .B(p_0_31[27]), .Cin(p_0_31[26]));
full_adder fa_1_31_2(.S(p_1_31[5]), .Cout(p_1_32[2]), .A(p_0_31[25]), .B(p_0_31[24]), .Cin(p_0_31[23]));
half_adder ha_1_31(.S(p_1_31[6]), .Cout(p_1_32[3]), .A(p_0_31[22]), .B(p_0_31[21]));
full_adder fa_1_32_0(.S(p_1_32[4]), .Cout(p_1_33[0]), .A(p_0_32[30]), .B(p_0_32[29]), .Cin(p_0_32[28]));
full_adder fa_1_32_1(.S(p_1_32[5]), .Cout(p_1_33[1]), .A(p_0_32[27]), .B(p_0_32[26]), .Cin(p_0_32[25]));
full_adder fa_1_32_2(.S(p_1_32[6]), .Cout(p_1_33[2]), .A(p_0_32[24]), .B(p_0_32[23]), .Cin(p_0_32[22]));
half_adder ha_1_32(.S(p_1_32[7]), .Cout(p_1_33[3]), .A(p_0_32[21]), .B(p_0_32[20]));
full_adder fa_1_33_0(.S(p_1_33[4]), .Cout(p_1_34[0]), .A(p_0_33[29]), .B(p_0_33[28]), .Cin(p_0_33[27]));
full_adder fa_1_33_1(.S(p_1_33[5]), .Cout(p_1_34[1]), .A(p_0_33[26]), .B(p_0_33[25]), .Cin(p_0_33[24]));
full_adder fa_1_33_2(.S(p_1_33[6]), .Cout(p_1_34[2]), .A(p_0_33[23]), .B(p_0_33[22]), .Cin(p_0_33[21]));
full_adder fa_1_34_0(.S(p_1_34[3]), .Cout(p_1_35[0]), .A(p_0_34[28]), .B(p_0_34[27]), .Cin(p_0_34[26]));
full_adder fa_1_34_1(.S(p_1_34[4]), .Cout(p_1_35[1]), .A(p_0_34[25]), .B(p_0_34[24]), .Cin(p_0_34[23]));
full_adder fa_1_35_0(.S(p_1_35[2]), .Cout(p_1_36[0]), .A(p_0_35[27]), .B(p_0_35[26]), .Cin(p_0_35[25]));

// Stage 2 non-added partial products
assign p_2_0[0:0] = p_1_0[0:0];
assign p_2_1[1:0] = p_1_1[1:0];
assign p_2_2[2:0] = p_1_2[2:0];
assign p_2_3[3:0] = p_1_3[3:0];
assign p_2_4[4:0] = p_1_4[4:0];
assign p_2_5[5:0] = p_1_5[5:0];
assign p_2_6[6:0] = p_1_6[6:0];
assign p_2_7[7:0] = p_1_7[7:0];
assign p_2_8[8:0] = p_1_8[8:0];
assign p_2_9[9:0] = p_1_9[9:0];
assign p_2_10[10:0] = p_1_10[10:0];
assign p_2_11[11:0] = p_1_11[11:0];
assign p_2_12[12:0] = p_1_12[12:0];
assign p_2_13[13:0] = p_1_13[13:0];
assign p_2_14[14:0] = p_1_14[14:0];
assign p_2_15[15:0] = p_1_15[15:0];
assign p_2_16[16:0] = p_1_16[16:0];
assign p_2_17[17:0] = p_1_17[17:0];
assign p_2_18[18:0] = p_1_18[18:0];
assign p_2_19[18:1] = p_1_19[17:0];
assign p_2_20[18:3] = p_1_20[15:0];
assign p_2_21[18:5] = p_1_21[13:0];
assign p_2_22[18:7] = p_1_22[11:0];
assign p_2_23[18:9] = p_1_23[9:0];
assign p_2_24[18:11] = p_1_24[7:0];
assign p_2_25[18:13] = p_1_25[5:0];
assign p_2_26[18:15] = p_1_26[3:0];
assign p_2_27[18:17] = p_1_27[1:0];
assign p_2_28[18:18] = p_1_28[0:0];
assign p_2_29[18:18] = p_1_29[0:0];
assign p_2_30[18:18] = p_1_30[0:0];
assign p_2_31[18:18] = p_1_31[0:0];
assign p_2_32[18:18] = p_1_32[0:0];
assign p_2_33[18:18] = p_1_33[0:0];
assign p_2_34[18:18] = p_1_34[0:0];
assign p_2_35[18:18] = p_1_35[0:0];
assign p_2_36[18:18] = p_1_36[0:0];
assign p_2_37[18:17] = p_1_37[1:0];
assign p_2_38[18:15] = p_1_38[3:0];
assign p_2_39[18:13] = p_1_39[5:0];
assign p_2_40[18:11] = p_1_40[7:0];
assign p_2_41[18:9] = p_1_41[9:0];
assign p_2_42[18:7] = p_1_42[11:0];
assign p_2_43[18:5] = p_1_43[13:0];
assign p_2_44[18:3] = p_1_44[15:0];
assign p_2_45[18:1] = p_1_45[17:0];
assign p_2_46[16:0] = p_1_46[16:0];
assign p_2_47[15:0] = p_1_47[15:0];
assign p_2_48[14:0] = p_1_48[14:0];
assign p_2_49[13:0] = p_1_49[13:0];
assign p_2_50[12:0] = p_1_50[12:0];
assign p_2_51[11:0] = p_1_51[11:0];
assign p_2_52[10:0] = p_1_52[10:0];
assign p_2_53[9:0] = p_1_53[9:0];
assign p_2_54[8:0] = p_1_54[8:0];
assign p_2_55[7:0] = p_1_55[7:0];
assign p_2_56[6:0] = p_1_56[6:0];
assign p_2_57[5:0] = p_1_57[5:0];
assign p_2_58[4:0] = p_1_58[4:0];
assign p_2_59[3:0] = p_1_59[3:0];
assign p_2_60[2:0] = p_1_60[2:0];
assign p_2_61[1:0] = p_1_61[1:0];
assign p_2_62[0:0] = p_1_62[0:0];
// Stage 2 adders
half_adder ha_2_19(.S(p_2_19[0]), .Cout(p_2_20[0]), .A(p_1_19[19]), .B(p_1_19[18]));
full_adder fa_2_20_0(.S(p_2_20[1]), .Cout(p_2_21[0]), .A(p_1_20[20]), .B(p_1_20[19]), .Cin(p_1_20[18]));
half_adder ha_2_20(.S(p_2_20[2]), .Cout(p_2_21[1]), .A(p_1_20[17]), .B(p_1_20[16]));
full_adder fa_2_21_0(.S(p_2_21[2]), .Cout(p_2_22[0]), .A(p_1_21[21]), .B(p_1_21[20]), .Cin(p_1_21[19]));
full_adder fa_2_21_1(.S(p_2_21[3]), .Cout(p_2_22[1]), .A(p_1_21[18]), .B(p_1_21[17]), .Cin(p_1_21[16]));
half_adder ha_2_21(.S(p_2_21[4]), .Cout(p_2_22[2]), .A(p_1_21[15]), .B(p_1_21[14]));
full_adder fa_2_22_0(.S(p_2_22[3]), .Cout(p_2_23[0]), .A(p_1_22[22]), .B(p_1_22[21]), .Cin(p_1_22[20]));
full_adder fa_2_22_1(.S(p_2_22[4]), .Cout(p_2_23[1]), .A(p_1_22[19]), .B(p_1_22[18]), .Cin(p_1_22[17]));
full_adder fa_2_22_2(.S(p_2_22[5]), .Cout(p_2_23[2]), .A(p_1_22[16]), .B(p_1_22[15]), .Cin(p_1_22[14]));
half_adder ha_2_22(.S(p_2_22[6]), .Cout(p_2_23[3]), .A(p_1_22[13]), .B(p_1_22[12]));
full_adder fa_2_23_0(.S(p_2_23[4]), .Cout(p_2_24[0]), .A(p_1_23[23]), .B(p_1_23[22]), .Cin(p_1_23[21]));
full_adder fa_2_23_1(.S(p_2_23[5]), .Cout(p_2_24[1]), .A(p_1_23[20]), .B(p_1_23[19]), .Cin(p_1_23[18]));
full_adder fa_2_23_2(.S(p_2_23[6]), .Cout(p_2_24[2]), .A(p_1_23[17]), .B(p_1_23[16]), .Cin(p_1_23[15]));
full_adder fa_2_23_3(.S(p_2_23[7]), .Cout(p_2_24[3]), .A(p_1_23[14]), .B(p_1_23[13]), .Cin(p_1_23[12]));
half_adder ha_2_23(.S(p_2_23[8]), .Cout(p_2_24[4]), .A(p_1_23[11]), .B(p_1_23[10]));
full_adder fa_2_24_0(.S(p_2_24[5]), .Cout(p_2_25[0]), .A(p_1_24[24]), .B(p_1_24[23]), .Cin(p_1_24[22]));
full_adder fa_2_24_1(.S(p_2_24[6]), .Cout(p_2_25[1]), .A(p_1_24[21]), .B(p_1_24[20]), .Cin(p_1_24[19]));
full_adder fa_2_24_2(.S(p_2_24[7]), .Cout(p_2_25[2]), .A(p_1_24[18]), .B(p_1_24[17]), .Cin(p_1_24[16]));
full_adder fa_2_24_3(.S(p_2_24[8]), .Cout(p_2_25[3]), .A(p_1_24[15]), .B(p_1_24[14]), .Cin(p_1_24[13]));
full_adder fa_2_24_4(.S(p_2_24[9]), .Cout(p_2_25[4]), .A(p_1_24[12]), .B(p_1_24[11]), .Cin(p_1_24[10]));
half_adder ha_2_24(.S(p_2_24[10]), .Cout(p_2_25[5]), .A(p_1_24[9]), .B(p_1_24[8]));
full_adder fa_2_25_0(.S(p_2_25[6]), .Cout(p_2_26[0]), .A(p_1_25[25]), .B(p_1_25[24]), .Cin(p_1_25[23]));
full_adder fa_2_25_1(.S(p_2_25[7]), .Cout(p_2_26[1]), .A(p_1_25[22]), .B(p_1_25[21]), .Cin(p_1_25[20]));
full_adder fa_2_25_2(.S(p_2_25[8]), .Cout(p_2_26[2]), .A(p_1_25[19]), .B(p_1_25[18]), .Cin(p_1_25[17]));
full_adder fa_2_25_3(.S(p_2_25[9]), .Cout(p_2_26[3]), .A(p_1_25[16]), .B(p_1_25[15]), .Cin(p_1_25[14]));
full_adder fa_2_25_4(.S(p_2_25[10]), .Cout(p_2_26[4]), .A(p_1_25[13]), .B(p_1_25[12]), .Cin(p_1_25[11]));
full_adder fa_2_25_5(.S(p_2_25[11]), .Cout(p_2_26[5]), .A(p_1_25[10]), .B(p_1_25[9]), .Cin(p_1_25[8]));
half_adder ha_2_25(.S(p_2_25[12]), .Cout(p_2_26[6]), .A(p_1_25[7]), .B(p_1_25[6]));
full_adder fa_2_26_0(.S(p_2_26[7]), .Cout(p_2_27[0]), .A(p_1_26[26]), .B(p_1_26[25]), .Cin(p_1_26[24]));
full_adder fa_2_26_1(.S(p_2_26[8]), .Cout(p_2_27[1]), .A(p_1_26[23]), .B(p_1_26[22]), .Cin(p_1_26[21]));
full_adder fa_2_26_2(.S(p_2_26[9]), .Cout(p_2_27[2]), .A(p_1_26[20]), .B(p_1_26[19]), .Cin(p_1_26[18]));
full_adder fa_2_26_3(.S(p_2_26[10]), .Cout(p_2_27[3]), .A(p_1_26[17]), .B(p_1_26[16]), .Cin(p_1_26[15]));
full_adder fa_2_26_4(.S(p_2_26[11]), .Cout(p_2_27[4]), .A(p_1_26[14]), .B(p_1_26[13]), .Cin(p_1_26[12]));
full_adder fa_2_26_5(.S(p_2_26[12]), .Cout(p_2_27[5]), .A(p_1_26[11]), .B(p_1_26[10]), .Cin(p_1_26[9]));
full_adder fa_2_26_6(.S(p_2_26[13]), .Cout(p_2_27[6]), .A(p_1_26[8]), .B(p_1_26[7]), .Cin(p_1_26[6]));
half_adder ha_2_26(.S(p_2_26[14]), .Cout(p_2_27[7]), .A(p_1_26[5]), .B(p_1_26[4]));
full_adder fa_2_27_0(.S(p_2_27[8]), .Cout(p_2_28[0]), .A(p_1_27[27]), .B(p_1_27[26]), .Cin(p_1_27[25]));
full_adder fa_2_27_1(.S(p_2_27[9]), .Cout(p_2_28[1]), .A(p_1_27[24]), .B(p_1_27[23]), .Cin(p_1_27[22]));
full_adder fa_2_27_2(.S(p_2_27[10]), .Cout(p_2_28[2]), .A(p_1_27[21]), .B(p_1_27[20]), .Cin(p_1_27[19]));
full_adder fa_2_27_3(.S(p_2_27[11]), .Cout(p_2_28[3]), .A(p_1_27[18]), .B(p_1_27[17]), .Cin(p_1_27[16]));
full_adder fa_2_27_4(.S(p_2_27[12]), .Cout(p_2_28[4]), .A(p_1_27[15]), .B(p_1_27[14]), .Cin(p_1_27[13]));
full_adder fa_2_27_5(.S(p_2_27[13]), .Cout(p_2_28[5]), .A(p_1_27[12]), .B(p_1_27[11]), .Cin(p_1_27[10]));
full_adder fa_2_27_6(.S(p_2_27[14]), .Cout(p_2_28[6]), .A(p_1_27[9]), .B(p_1_27[8]), .Cin(p_1_27[7]));
full_adder fa_2_27_7(.S(p_2_27[15]), .Cout(p_2_28[7]), .A(p_1_27[6]), .B(p_1_27[5]), .Cin(p_1_27[4]));
half_adder ha_2_27(.S(p_2_27[16]), .Cout(p_2_28[8]), .A(p_1_27[3]), .B(p_1_27[2]));
full_adder fa_2_28_0(.S(p_2_28[9]), .Cout(p_2_29[0]), .A(p_1_28[27]), .B(p_1_28[26]), .Cin(p_1_28[25]));
full_adder fa_2_28_1(.S(p_2_28[10]), .Cout(p_2_29[1]), .A(p_1_28[24]), .B(p_1_28[23]), .Cin(p_1_28[22]));
full_adder fa_2_28_2(.S(p_2_28[11]), .Cout(p_2_29[2]), .A(p_1_28[21]), .B(p_1_28[20]), .Cin(p_1_28[19]));
full_adder fa_2_28_3(.S(p_2_28[12]), .Cout(p_2_29[3]), .A(p_1_28[18]), .B(p_1_28[17]), .Cin(p_1_28[16]));
full_adder fa_2_28_4(.S(p_2_28[13]), .Cout(p_2_29[4]), .A(p_1_28[15]), .B(p_1_28[14]), .Cin(p_1_28[13]));
full_adder fa_2_28_5(.S(p_2_28[14]), .Cout(p_2_29[5]), .A(p_1_28[12]), .B(p_1_28[11]), .Cin(p_1_28[10]));
full_adder fa_2_28_6(.S(p_2_28[15]), .Cout(p_2_29[6]), .A(p_1_28[9]), .B(p_1_28[8]), .Cin(p_1_28[7]));
full_adder fa_2_28_7(.S(p_2_28[16]), .Cout(p_2_29[7]), .A(p_1_28[6]), .B(p_1_28[5]), .Cin(p_1_28[4]));
full_adder fa_2_28_8(.S(p_2_28[17]), .Cout(p_2_29[8]), .A(p_1_28[3]), .B(p_1_28[2]), .Cin(p_1_28[1]));
full_adder fa_2_29_0(.S(p_2_29[9]), .Cout(p_2_30[0]), .A(p_1_29[27]), .B(p_1_29[26]), .Cin(p_1_29[25]));
full_adder fa_2_29_1(.S(p_2_29[10]), .Cout(p_2_30[1]), .A(p_1_29[24]), .B(p_1_29[23]), .Cin(p_1_29[22]));
full_adder fa_2_29_2(.S(p_2_29[11]), .Cout(p_2_30[2]), .A(p_1_29[21]), .B(p_1_29[20]), .Cin(p_1_29[19]));
full_adder fa_2_29_3(.S(p_2_29[12]), .Cout(p_2_30[3]), .A(p_1_29[18]), .B(p_1_29[17]), .Cin(p_1_29[16]));
full_adder fa_2_29_4(.S(p_2_29[13]), .Cout(p_2_30[4]), .A(p_1_29[15]), .B(p_1_29[14]), .Cin(p_1_29[13]));
full_adder fa_2_29_5(.S(p_2_29[14]), .Cout(p_2_30[5]), .A(p_1_29[12]), .B(p_1_29[11]), .Cin(p_1_29[10]));
full_adder fa_2_29_6(.S(p_2_29[15]), .Cout(p_2_30[6]), .A(p_1_29[9]), .B(p_1_29[8]), .Cin(p_1_29[7]));
full_adder fa_2_29_7(.S(p_2_29[16]), .Cout(p_2_30[7]), .A(p_1_29[6]), .B(p_1_29[5]), .Cin(p_1_29[4]));
full_adder fa_2_29_8(.S(p_2_29[17]), .Cout(p_2_30[8]), .A(p_1_29[3]), .B(p_1_29[2]), .Cin(p_1_29[1]));
full_adder fa_2_30_0(.S(p_2_30[9]), .Cout(p_2_31[0]), .A(p_1_30[27]), .B(p_1_30[26]), .Cin(p_1_30[25]));
full_adder fa_2_30_1(.S(p_2_30[10]), .Cout(p_2_31[1]), .A(p_1_30[24]), .B(p_1_30[23]), .Cin(p_1_30[22]));
full_adder fa_2_30_2(.S(p_2_30[11]), .Cout(p_2_31[2]), .A(p_1_30[21]), .B(p_1_30[20]), .Cin(p_1_30[19]));
full_adder fa_2_30_3(.S(p_2_30[12]), .Cout(p_2_31[3]), .A(p_1_30[18]), .B(p_1_30[17]), .Cin(p_1_30[16]));
full_adder fa_2_30_4(.S(p_2_30[13]), .Cout(p_2_31[4]), .A(p_1_30[15]), .B(p_1_30[14]), .Cin(p_1_30[13]));
full_adder fa_2_30_5(.S(p_2_30[14]), .Cout(p_2_31[5]), .A(p_1_30[12]), .B(p_1_30[11]), .Cin(p_1_30[10]));
full_adder fa_2_30_6(.S(p_2_30[15]), .Cout(p_2_31[6]), .A(p_1_30[9]), .B(p_1_30[8]), .Cin(p_1_30[7]));
full_adder fa_2_30_7(.S(p_2_30[16]), .Cout(p_2_31[7]), .A(p_1_30[6]), .B(p_1_30[5]), .Cin(p_1_30[4]));
full_adder fa_2_30_8(.S(p_2_30[17]), .Cout(p_2_31[8]), .A(p_1_30[3]), .B(p_1_30[2]), .Cin(p_1_30[1]));
full_adder fa_2_31_0(.S(p_2_31[9]), .Cout(p_2_32[0]), .A(p_1_31[27]), .B(p_1_31[26]), .Cin(p_1_31[25]));
full_adder fa_2_31_1(.S(p_2_31[10]), .Cout(p_2_32[1]), .A(p_1_31[24]), .B(p_1_31[23]), .Cin(p_1_31[22]));
full_adder fa_2_31_2(.S(p_2_31[11]), .Cout(p_2_32[2]), .A(p_1_31[21]), .B(p_1_31[20]), .Cin(p_1_31[19]));
full_adder fa_2_31_3(.S(p_2_31[12]), .Cout(p_2_32[3]), .A(p_1_31[18]), .B(p_1_31[17]), .Cin(p_1_31[16]));
full_adder fa_2_31_4(.S(p_2_31[13]), .Cout(p_2_32[4]), .A(p_1_31[15]), .B(p_1_31[14]), .Cin(p_1_31[13]));
full_adder fa_2_31_5(.S(p_2_31[14]), .Cout(p_2_32[5]), .A(p_1_31[12]), .B(p_1_31[11]), .Cin(p_1_31[10]));
full_adder fa_2_31_6(.S(p_2_31[15]), .Cout(p_2_32[6]), .A(p_1_31[9]), .B(p_1_31[8]), .Cin(p_1_31[7]));
full_adder fa_2_31_7(.S(p_2_31[16]), .Cout(p_2_32[7]), .A(p_1_31[6]), .B(p_1_31[5]), .Cin(p_1_31[4]));
full_adder fa_2_31_8(.S(p_2_31[17]), .Cout(p_2_32[8]), .A(p_1_31[3]), .B(p_1_31[2]), .Cin(p_1_31[1]));
full_adder fa_2_32_0(.S(p_2_32[9]), .Cout(p_2_33[0]), .A(p_1_32[27]), .B(p_1_32[26]), .Cin(p_1_32[25]));
full_adder fa_2_32_1(.S(p_2_32[10]), .Cout(p_2_33[1]), .A(p_1_32[24]), .B(p_1_32[23]), .Cin(p_1_32[22]));
full_adder fa_2_32_2(.S(p_2_32[11]), .Cout(p_2_33[2]), .A(p_1_32[21]), .B(p_1_32[20]), .Cin(p_1_32[19]));
full_adder fa_2_32_3(.S(p_2_32[12]), .Cout(p_2_33[3]), .A(p_1_32[18]), .B(p_1_32[17]), .Cin(p_1_32[16]));
full_adder fa_2_32_4(.S(p_2_32[13]), .Cout(p_2_33[4]), .A(p_1_32[15]), .B(p_1_32[14]), .Cin(p_1_32[13]));
full_adder fa_2_32_5(.S(p_2_32[14]), .Cout(p_2_33[5]), .A(p_1_32[12]), .B(p_1_32[11]), .Cin(p_1_32[10]));
full_adder fa_2_32_6(.S(p_2_32[15]), .Cout(p_2_33[6]), .A(p_1_32[9]), .B(p_1_32[8]), .Cin(p_1_32[7]));
full_adder fa_2_32_7(.S(p_2_32[16]), .Cout(p_2_33[7]), .A(p_1_32[6]), .B(p_1_32[5]), .Cin(p_1_32[4]));
full_adder fa_2_32_8(.S(p_2_32[17]), .Cout(p_2_33[8]), .A(p_1_32[3]), .B(p_1_32[2]), .Cin(p_1_32[1]));
full_adder fa_2_33_0(.S(p_2_33[9]), .Cout(p_2_34[0]), .A(p_1_33[27]), .B(p_1_33[26]), .Cin(p_1_33[25]));
full_adder fa_2_33_1(.S(p_2_33[10]), .Cout(p_2_34[1]), .A(p_1_33[24]), .B(p_1_33[23]), .Cin(p_1_33[22]));
full_adder fa_2_33_2(.S(p_2_33[11]), .Cout(p_2_34[2]), .A(p_1_33[21]), .B(p_1_33[20]), .Cin(p_1_33[19]));
full_adder fa_2_33_3(.S(p_2_33[12]), .Cout(p_2_34[3]), .A(p_1_33[18]), .B(p_1_33[17]), .Cin(p_1_33[16]));
full_adder fa_2_33_4(.S(p_2_33[13]), .Cout(p_2_34[4]), .A(p_1_33[15]), .B(p_1_33[14]), .Cin(p_1_33[13]));
full_adder fa_2_33_5(.S(p_2_33[14]), .Cout(p_2_34[5]), .A(p_1_33[12]), .B(p_1_33[11]), .Cin(p_1_33[10]));
full_adder fa_2_33_6(.S(p_2_33[15]), .Cout(p_2_34[6]), .A(p_1_33[9]), .B(p_1_33[8]), .Cin(p_1_33[7]));
full_adder fa_2_33_7(.S(p_2_33[16]), .Cout(p_2_34[7]), .A(p_1_33[6]), .B(p_1_33[5]), .Cin(p_1_33[4]));
full_adder fa_2_33_8(.S(p_2_33[17]), .Cout(p_2_34[8]), .A(p_1_33[3]), .B(p_1_33[2]), .Cin(p_1_33[1]));
full_adder fa_2_34_0(.S(p_2_34[9]), .Cout(p_2_35[0]), .A(p_1_34[27]), .B(p_1_34[26]), .Cin(p_1_34[25]));
full_adder fa_2_34_1(.S(p_2_34[10]), .Cout(p_2_35[1]), .A(p_1_34[24]), .B(p_1_34[23]), .Cin(p_1_34[22]));
full_adder fa_2_34_2(.S(p_2_34[11]), .Cout(p_2_35[2]), .A(p_1_34[21]), .B(p_1_34[20]), .Cin(p_1_34[19]));
full_adder fa_2_34_3(.S(p_2_34[12]), .Cout(p_2_35[3]), .A(p_1_34[18]), .B(p_1_34[17]), .Cin(p_1_34[16]));
full_adder fa_2_34_4(.S(p_2_34[13]), .Cout(p_2_35[4]), .A(p_1_34[15]), .B(p_1_34[14]), .Cin(p_1_34[13]));
full_adder fa_2_34_5(.S(p_2_34[14]), .Cout(p_2_35[5]), .A(p_1_34[12]), .B(p_1_34[11]), .Cin(p_1_34[10]));
full_adder fa_2_34_6(.S(p_2_34[15]), .Cout(p_2_35[6]), .A(p_1_34[9]), .B(p_1_34[8]), .Cin(p_1_34[7]));
full_adder fa_2_34_7(.S(p_2_34[16]), .Cout(p_2_35[7]), .A(p_1_34[6]), .B(p_1_34[5]), .Cin(p_1_34[4]));
full_adder fa_2_34_8(.S(p_2_34[17]), .Cout(p_2_35[8]), .A(p_1_34[3]), .B(p_1_34[2]), .Cin(p_1_34[1]));
full_adder fa_2_35_0(.S(p_2_35[9]), .Cout(p_2_36[0]), .A(p_1_35[27]), .B(p_1_35[26]), .Cin(p_1_35[25]));
full_adder fa_2_35_1(.S(p_2_35[10]), .Cout(p_2_36[1]), .A(p_1_35[24]), .B(p_1_35[23]), .Cin(p_1_35[22]));
full_adder fa_2_35_2(.S(p_2_35[11]), .Cout(p_2_36[2]), .A(p_1_35[21]), .B(p_1_35[20]), .Cin(p_1_35[19]));
full_adder fa_2_35_3(.S(p_2_35[12]), .Cout(p_2_36[3]), .A(p_1_35[18]), .B(p_1_35[17]), .Cin(p_1_35[16]));
full_adder fa_2_35_4(.S(p_2_35[13]), .Cout(p_2_36[4]), .A(p_1_35[15]), .B(p_1_35[14]), .Cin(p_1_35[13]));
full_adder fa_2_35_5(.S(p_2_35[14]), .Cout(p_2_36[5]), .A(p_1_35[12]), .B(p_1_35[11]), .Cin(p_1_35[10]));
full_adder fa_2_35_6(.S(p_2_35[15]), .Cout(p_2_36[6]), .A(p_1_35[9]), .B(p_1_35[8]), .Cin(p_1_35[7]));
full_adder fa_2_35_7(.S(p_2_35[16]), .Cout(p_2_36[7]), .A(p_1_35[6]), .B(p_1_35[5]), .Cin(p_1_35[4]));
full_adder fa_2_35_8(.S(p_2_35[17]), .Cout(p_2_36[8]), .A(p_1_35[3]), .B(p_1_35[2]), .Cin(p_1_35[1]));
full_adder fa_2_36_0(.S(p_2_36[9]), .Cout(p_2_37[0]), .A(p_1_36[27]), .B(p_1_36[26]), .Cin(p_1_36[25]));
full_adder fa_2_36_1(.S(p_2_36[10]), .Cout(p_2_37[1]), .A(p_1_36[24]), .B(p_1_36[23]), .Cin(p_1_36[22]));
full_adder fa_2_36_2(.S(p_2_36[11]), .Cout(p_2_37[2]), .A(p_1_36[21]), .B(p_1_36[20]), .Cin(p_1_36[19]));
full_adder fa_2_36_3(.S(p_2_36[12]), .Cout(p_2_37[3]), .A(p_1_36[18]), .B(p_1_36[17]), .Cin(p_1_36[16]));
full_adder fa_2_36_4(.S(p_2_36[13]), .Cout(p_2_37[4]), .A(p_1_36[15]), .B(p_1_36[14]), .Cin(p_1_36[13]));
full_adder fa_2_36_5(.S(p_2_36[14]), .Cout(p_2_37[5]), .A(p_1_36[12]), .B(p_1_36[11]), .Cin(p_1_36[10]));
full_adder fa_2_36_6(.S(p_2_36[15]), .Cout(p_2_37[6]), .A(p_1_36[9]), .B(p_1_36[8]), .Cin(p_1_36[7]));
full_adder fa_2_36_7(.S(p_2_36[16]), .Cout(p_2_37[7]), .A(p_1_36[6]), .B(p_1_36[5]), .Cin(p_1_36[4]));
full_adder fa_2_36_8(.S(p_2_36[17]), .Cout(p_2_37[8]), .A(p_1_36[3]), .B(p_1_36[2]), .Cin(p_1_36[1]));
full_adder fa_2_37_0(.S(p_2_37[9]), .Cout(p_2_38[0]), .A(p_1_37[25]), .B(p_1_37[24]), .Cin(p_1_37[23]));
full_adder fa_2_37_1(.S(p_2_37[10]), .Cout(p_2_38[1]), .A(p_1_37[22]), .B(p_1_37[21]), .Cin(p_1_37[20]));
full_adder fa_2_37_2(.S(p_2_37[11]), .Cout(p_2_38[2]), .A(p_1_37[19]), .B(p_1_37[18]), .Cin(p_1_37[17]));
full_adder fa_2_37_3(.S(p_2_37[12]), .Cout(p_2_38[3]), .A(p_1_37[16]), .B(p_1_37[15]), .Cin(p_1_37[14]));
full_adder fa_2_37_4(.S(p_2_37[13]), .Cout(p_2_38[4]), .A(p_1_37[13]), .B(p_1_37[12]), .Cin(p_1_37[11]));
full_adder fa_2_37_5(.S(p_2_37[14]), .Cout(p_2_38[5]), .A(p_1_37[10]), .B(p_1_37[9]), .Cin(p_1_37[8]));
full_adder fa_2_37_6(.S(p_2_37[15]), .Cout(p_2_38[6]), .A(p_1_37[7]), .B(p_1_37[6]), .Cin(p_1_37[5]));
full_adder fa_2_37_7(.S(p_2_37[16]), .Cout(p_2_38[7]), .A(p_1_37[4]), .B(p_1_37[3]), .Cin(p_1_37[2]));
full_adder fa_2_38_0(.S(p_2_38[8]), .Cout(p_2_39[0]), .A(p_1_38[24]), .B(p_1_38[23]), .Cin(p_1_38[22]));
full_adder fa_2_38_1(.S(p_2_38[9]), .Cout(p_2_39[1]), .A(p_1_38[21]), .B(p_1_38[20]), .Cin(p_1_38[19]));
full_adder fa_2_38_2(.S(p_2_38[10]), .Cout(p_2_39[2]), .A(p_1_38[18]), .B(p_1_38[17]), .Cin(p_1_38[16]));
full_adder fa_2_38_3(.S(p_2_38[11]), .Cout(p_2_39[3]), .A(p_1_38[15]), .B(p_1_38[14]), .Cin(p_1_38[13]));
full_adder fa_2_38_4(.S(p_2_38[12]), .Cout(p_2_39[4]), .A(p_1_38[12]), .B(p_1_38[11]), .Cin(p_1_38[10]));
full_adder fa_2_38_5(.S(p_2_38[13]), .Cout(p_2_39[5]), .A(p_1_38[9]), .B(p_1_38[8]), .Cin(p_1_38[7]));
full_adder fa_2_38_6(.S(p_2_38[14]), .Cout(p_2_39[6]), .A(p_1_38[6]), .B(p_1_38[5]), .Cin(p_1_38[4]));
full_adder fa_2_39_0(.S(p_2_39[7]), .Cout(p_2_40[0]), .A(p_1_39[23]), .B(p_1_39[22]), .Cin(p_1_39[21]));
full_adder fa_2_39_1(.S(p_2_39[8]), .Cout(p_2_40[1]), .A(p_1_39[20]), .B(p_1_39[19]), .Cin(p_1_39[18]));
full_adder fa_2_39_2(.S(p_2_39[9]), .Cout(p_2_40[2]), .A(p_1_39[17]), .B(p_1_39[16]), .Cin(p_1_39[15]));
full_adder fa_2_39_3(.S(p_2_39[10]), .Cout(p_2_40[3]), .A(p_1_39[14]), .B(p_1_39[13]), .Cin(p_1_39[12]));
full_adder fa_2_39_4(.S(p_2_39[11]), .Cout(p_2_40[4]), .A(p_1_39[11]), .B(p_1_39[10]), .Cin(p_1_39[9]));
full_adder fa_2_39_5(.S(p_2_39[12]), .Cout(p_2_40[5]), .A(p_1_39[8]), .B(p_1_39[7]), .Cin(p_1_39[6]));
full_adder fa_2_40_0(.S(p_2_40[6]), .Cout(p_2_41[0]), .A(p_1_40[22]), .B(p_1_40[21]), .Cin(p_1_40[20]));
full_adder fa_2_40_1(.S(p_2_40[7]), .Cout(p_2_41[1]), .A(p_1_40[19]), .B(p_1_40[18]), .Cin(p_1_40[17]));
full_adder fa_2_40_2(.S(p_2_40[8]), .Cout(p_2_41[2]), .A(p_1_40[16]), .B(p_1_40[15]), .Cin(p_1_40[14]));
full_adder fa_2_40_3(.S(p_2_40[9]), .Cout(p_2_41[3]), .A(p_1_40[13]), .B(p_1_40[12]), .Cin(p_1_40[11]));
full_adder fa_2_40_4(.S(p_2_40[10]), .Cout(p_2_41[4]), .A(p_1_40[10]), .B(p_1_40[9]), .Cin(p_1_40[8]));
full_adder fa_2_41_0(.S(p_2_41[5]), .Cout(p_2_42[0]), .A(p_1_41[21]), .B(p_1_41[20]), .Cin(p_1_41[19]));
full_adder fa_2_41_1(.S(p_2_41[6]), .Cout(p_2_42[1]), .A(p_1_41[18]), .B(p_1_41[17]), .Cin(p_1_41[16]));
full_adder fa_2_41_2(.S(p_2_41[7]), .Cout(p_2_42[2]), .A(p_1_41[15]), .B(p_1_41[14]), .Cin(p_1_41[13]));
full_adder fa_2_41_3(.S(p_2_41[8]), .Cout(p_2_42[3]), .A(p_1_41[12]), .B(p_1_41[11]), .Cin(p_1_41[10]));
full_adder fa_2_42_0(.S(p_2_42[4]), .Cout(p_2_43[0]), .A(p_1_42[20]), .B(p_1_42[19]), .Cin(p_1_42[18]));
full_adder fa_2_42_1(.S(p_2_42[5]), .Cout(p_2_43[1]), .A(p_1_42[17]), .B(p_1_42[16]), .Cin(p_1_42[15]));
full_adder fa_2_42_2(.S(p_2_42[6]), .Cout(p_2_43[2]), .A(p_1_42[14]), .B(p_1_42[13]), .Cin(p_1_42[12]));
full_adder fa_2_43_0(.S(p_2_43[3]), .Cout(p_2_44[0]), .A(p_1_43[19]), .B(p_1_43[18]), .Cin(p_1_43[17]));
full_adder fa_2_43_1(.S(p_2_43[4]), .Cout(p_2_44[1]), .A(p_1_43[16]), .B(p_1_43[15]), .Cin(p_1_43[14]));
full_adder fa_2_44_0(.S(p_2_44[2]), .Cout(p_2_45[0]), .A(p_1_44[18]), .B(p_1_44[17]), .Cin(p_1_44[16]));

// Stage 3 non-added partial products
assign p_3_0[0:0] = p_2_0[0:0];
assign p_3_1[1:0] = p_2_1[1:0];
assign p_3_2[2:0] = p_2_2[2:0];
assign p_3_3[3:0] = p_2_3[3:0];
assign p_3_4[4:0] = p_2_4[4:0];
assign p_3_5[5:0] = p_2_5[5:0];
assign p_3_6[6:0] = p_2_6[6:0];
assign p_3_7[7:0] = p_2_7[7:0];
assign p_3_8[8:0] = p_2_8[8:0];
assign p_3_9[9:0] = p_2_9[9:0];
assign p_3_10[10:0] = p_2_10[10:0];
assign p_3_11[11:0] = p_2_11[11:0];
assign p_3_12[12:0] = p_2_12[12:0];
assign p_3_13[12:1] = p_2_13[11:0];
assign p_3_14[12:3] = p_2_14[9:0];
assign p_3_15[12:5] = p_2_15[7:0];
assign p_3_16[12:7] = p_2_16[5:0];
assign p_3_17[12:9] = p_2_17[3:0];
assign p_3_18[12:11] = p_2_18[1:0];
assign p_3_19[12:12] = p_2_19[0:0];
assign p_3_20[12:12] = p_2_20[0:0];
assign p_3_21[12:12] = p_2_21[0:0];
assign p_3_22[12:12] = p_2_22[0:0];
assign p_3_23[12:12] = p_2_23[0:0];
assign p_3_24[12:12] = p_2_24[0:0];
assign p_3_25[12:12] = p_2_25[0:0];
assign p_3_26[12:12] = p_2_26[0:0];
assign p_3_27[12:12] = p_2_27[0:0];
assign p_3_28[12:12] = p_2_28[0:0];
assign p_3_29[12:12] = p_2_29[0:0];
assign p_3_30[12:12] = p_2_30[0:0];
assign p_3_31[12:12] = p_2_31[0:0];
assign p_3_32[12:12] = p_2_32[0:0];
assign p_3_33[12:12] = p_2_33[0:0];
assign p_3_34[12:12] = p_2_34[0:0];
assign p_3_35[12:12] = p_2_35[0:0];
assign p_3_36[12:12] = p_2_36[0:0];
assign p_3_37[12:12] = p_2_37[0:0];
assign p_3_38[12:12] = p_2_38[0:0];
assign p_3_39[12:12] = p_2_39[0:0];
assign p_3_40[12:12] = p_2_40[0:0];
assign p_3_41[12:12] = p_2_41[0:0];
assign p_3_42[12:12] = p_2_42[0:0];
assign p_3_43[12:12] = p_2_43[0:0];
assign p_3_44[12:12] = p_2_44[0:0];
assign p_3_45[12:12] = p_2_45[0:0];
assign p_3_46[12:11] = p_2_46[1:0];
assign p_3_47[12:9] = p_2_47[3:0];
assign p_3_48[12:7] = p_2_48[5:0];
assign p_3_49[12:5] = p_2_49[7:0];
assign p_3_50[12:3] = p_2_50[9:0];
assign p_3_51[12:1] = p_2_51[11:0];
assign p_3_52[10:0] = p_2_52[10:0];
assign p_3_53[9:0] = p_2_53[9:0];
assign p_3_54[8:0] = p_2_54[8:0];
assign p_3_55[7:0] = p_2_55[7:0];
assign p_3_56[6:0] = p_2_56[6:0];
assign p_3_57[5:0] = p_2_57[5:0];
assign p_3_58[4:0] = p_2_58[4:0];
assign p_3_59[3:0] = p_2_59[3:0];
assign p_3_60[2:0] = p_2_60[2:0];
assign p_3_61[1:0] = p_2_61[1:0];
assign p_3_62[0:0] = p_2_62[0:0];
// Stage 3 adders
half_adder ha_3_13(.S(p_3_13[0]), .Cout(p_3_14[0]), .A(p_2_13[13]), .B(p_2_13[12]));
full_adder fa_3_14_0(.S(p_3_14[1]), .Cout(p_3_15[0]), .A(p_2_14[14]), .B(p_2_14[13]), .Cin(p_2_14[12]));
half_adder ha_3_14(.S(p_3_14[2]), .Cout(p_3_15[1]), .A(p_2_14[11]), .B(p_2_14[10]));
full_adder fa_3_15_0(.S(p_3_15[2]), .Cout(p_3_16[0]), .A(p_2_15[15]), .B(p_2_15[14]), .Cin(p_2_15[13]));
full_adder fa_3_15_1(.S(p_3_15[3]), .Cout(p_3_16[1]), .A(p_2_15[12]), .B(p_2_15[11]), .Cin(p_2_15[10]));
half_adder ha_3_15(.S(p_3_15[4]), .Cout(p_3_16[2]), .A(p_2_15[9]), .B(p_2_15[8]));
full_adder fa_3_16_0(.S(p_3_16[3]), .Cout(p_3_17[0]), .A(p_2_16[16]), .B(p_2_16[15]), .Cin(p_2_16[14]));
full_adder fa_3_16_1(.S(p_3_16[4]), .Cout(p_3_17[1]), .A(p_2_16[13]), .B(p_2_16[12]), .Cin(p_2_16[11]));
full_adder fa_3_16_2(.S(p_3_16[5]), .Cout(p_3_17[2]), .A(p_2_16[10]), .B(p_2_16[9]), .Cin(p_2_16[8]));
half_adder ha_3_16(.S(p_3_16[6]), .Cout(p_3_17[3]), .A(p_2_16[7]), .B(p_2_16[6]));
full_adder fa_3_17_0(.S(p_3_17[4]), .Cout(p_3_18[0]), .A(p_2_17[17]), .B(p_2_17[16]), .Cin(p_2_17[15]));
full_adder fa_3_17_1(.S(p_3_17[5]), .Cout(p_3_18[1]), .A(p_2_17[14]), .B(p_2_17[13]), .Cin(p_2_17[12]));
full_adder fa_3_17_2(.S(p_3_17[6]), .Cout(p_3_18[2]), .A(p_2_17[11]), .B(p_2_17[10]), .Cin(p_2_17[9]));
full_adder fa_3_17_3(.S(p_3_17[7]), .Cout(p_3_18[3]), .A(p_2_17[8]), .B(p_2_17[7]), .Cin(p_2_17[6]));
half_adder ha_3_17(.S(p_3_17[8]), .Cout(p_3_18[4]), .A(p_2_17[5]), .B(p_2_17[4]));
full_adder fa_3_18_0(.S(p_3_18[5]), .Cout(p_3_19[0]), .A(p_2_18[18]), .B(p_2_18[17]), .Cin(p_2_18[16]));
full_adder fa_3_18_1(.S(p_3_18[6]), .Cout(p_3_19[1]), .A(p_2_18[15]), .B(p_2_18[14]), .Cin(p_2_18[13]));
full_adder fa_3_18_2(.S(p_3_18[7]), .Cout(p_3_19[2]), .A(p_2_18[12]), .B(p_2_18[11]), .Cin(p_2_18[10]));
full_adder fa_3_18_3(.S(p_3_18[8]), .Cout(p_3_19[3]), .A(p_2_18[9]), .B(p_2_18[8]), .Cin(p_2_18[7]));
full_adder fa_3_18_4(.S(p_3_18[9]), .Cout(p_3_19[4]), .A(p_2_18[6]), .B(p_2_18[5]), .Cin(p_2_18[4]));
half_adder ha_3_18(.S(p_3_18[10]), .Cout(p_3_19[5]), .A(p_2_18[3]), .B(p_2_18[2]));
full_adder fa_3_19_0(.S(p_3_19[6]), .Cout(p_3_20[0]), .A(p_2_19[18]), .B(p_2_19[17]), .Cin(p_2_19[16]));
full_adder fa_3_19_1(.S(p_3_19[7]), .Cout(p_3_20[1]), .A(p_2_19[15]), .B(p_2_19[14]), .Cin(p_2_19[13]));
full_adder fa_3_19_2(.S(p_3_19[8]), .Cout(p_3_20[2]), .A(p_2_19[12]), .B(p_2_19[11]), .Cin(p_2_19[10]));
full_adder fa_3_19_3(.S(p_3_19[9]), .Cout(p_3_20[3]), .A(p_2_19[9]), .B(p_2_19[8]), .Cin(p_2_19[7]));
full_adder fa_3_19_4(.S(p_3_19[10]), .Cout(p_3_20[4]), .A(p_2_19[6]), .B(p_2_19[5]), .Cin(p_2_19[4]));
full_adder fa_3_19_5(.S(p_3_19[11]), .Cout(p_3_20[5]), .A(p_2_19[3]), .B(p_2_19[2]), .Cin(p_2_19[1]));
full_adder fa_3_20_0(.S(p_3_20[6]), .Cout(p_3_21[0]), .A(p_2_20[18]), .B(p_2_20[17]), .Cin(p_2_20[16]));
full_adder fa_3_20_1(.S(p_3_20[7]), .Cout(p_3_21[1]), .A(p_2_20[15]), .B(p_2_20[14]), .Cin(p_2_20[13]));
full_adder fa_3_20_2(.S(p_3_20[8]), .Cout(p_3_21[2]), .A(p_2_20[12]), .B(p_2_20[11]), .Cin(p_2_20[10]));
full_adder fa_3_20_3(.S(p_3_20[9]), .Cout(p_3_21[3]), .A(p_2_20[9]), .B(p_2_20[8]), .Cin(p_2_20[7]));
full_adder fa_3_20_4(.S(p_3_20[10]), .Cout(p_3_21[4]), .A(p_2_20[6]), .B(p_2_20[5]), .Cin(p_2_20[4]));
full_adder fa_3_20_5(.S(p_3_20[11]), .Cout(p_3_21[5]), .A(p_2_20[3]), .B(p_2_20[2]), .Cin(p_2_20[1]));
full_adder fa_3_21_0(.S(p_3_21[6]), .Cout(p_3_22[0]), .A(p_2_21[18]), .B(p_2_21[17]), .Cin(p_2_21[16]));
full_adder fa_3_21_1(.S(p_3_21[7]), .Cout(p_3_22[1]), .A(p_2_21[15]), .B(p_2_21[14]), .Cin(p_2_21[13]));
full_adder fa_3_21_2(.S(p_3_21[8]), .Cout(p_3_22[2]), .A(p_2_21[12]), .B(p_2_21[11]), .Cin(p_2_21[10]));
full_adder fa_3_21_3(.S(p_3_21[9]), .Cout(p_3_22[3]), .A(p_2_21[9]), .B(p_2_21[8]), .Cin(p_2_21[7]));
full_adder fa_3_21_4(.S(p_3_21[10]), .Cout(p_3_22[4]), .A(p_2_21[6]), .B(p_2_21[5]), .Cin(p_2_21[4]));
full_adder fa_3_21_5(.S(p_3_21[11]), .Cout(p_3_22[5]), .A(p_2_21[3]), .B(p_2_21[2]), .Cin(p_2_21[1]));
full_adder fa_3_22_0(.S(p_3_22[6]), .Cout(p_3_23[0]), .A(p_2_22[18]), .B(p_2_22[17]), .Cin(p_2_22[16]));
full_adder fa_3_22_1(.S(p_3_22[7]), .Cout(p_3_23[1]), .A(p_2_22[15]), .B(p_2_22[14]), .Cin(p_2_22[13]));
full_adder fa_3_22_2(.S(p_3_22[8]), .Cout(p_3_23[2]), .A(p_2_22[12]), .B(p_2_22[11]), .Cin(p_2_22[10]));
full_adder fa_3_22_3(.S(p_3_22[9]), .Cout(p_3_23[3]), .A(p_2_22[9]), .B(p_2_22[8]), .Cin(p_2_22[7]));
full_adder fa_3_22_4(.S(p_3_22[10]), .Cout(p_3_23[4]), .A(p_2_22[6]), .B(p_2_22[5]), .Cin(p_2_22[4]));
full_adder fa_3_22_5(.S(p_3_22[11]), .Cout(p_3_23[5]), .A(p_2_22[3]), .B(p_2_22[2]), .Cin(p_2_22[1]));
full_adder fa_3_23_0(.S(p_3_23[6]), .Cout(p_3_24[0]), .A(p_2_23[18]), .B(p_2_23[17]), .Cin(p_2_23[16]));
full_adder fa_3_23_1(.S(p_3_23[7]), .Cout(p_3_24[1]), .A(p_2_23[15]), .B(p_2_23[14]), .Cin(p_2_23[13]));
full_adder fa_3_23_2(.S(p_3_23[8]), .Cout(p_3_24[2]), .A(p_2_23[12]), .B(p_2_23[11]), .Cin(p_2_23[10]));
full_adder fa_3_23_3(.S(p_3_23[9]), .Cout(p_3_24[3]), .A(p_2_23[9]), .B(p_2_23[8]), .Cin(p_2_23[7]));
full_adder fa_3_23_4(.S(p_3_23[10]), .Cout(p_3_24[4]), .A(p_2_23[6]), .B(p_2_23[5]), .Cin(p_2_23[4]));
full_adder fa_3_23_5(.S(p_3_23[11]), .Cout(p_3_24[5]), .A(p_2_23[3]), .B(p_2_23[2]), .Cin(p_2_23[1]));
full_adder fa_3_24_0(.S(p_3_24[6]), .Cout(p_3_25[0]), .A(p_2_24[18]), .B(p_2_24[17]), .Cin(p_2_24[16]));
full_adder fa_3_24_1(.S(p_3_24[7]), .Cout(p_3_25[1]), .A(p_2_24[15]), .B(p_2_24[14]), .Cin(p_2_24[13]));
full_adder fa_3_24_2(.S(p_3_24[8]), .Cout(p_3_25[2]), .A(p_2_24[12]), .B(p_2_24[11]), .Cin(p_2_24[10]));
full_adder fa_3_24_3(.S(p_3_24[9]), .Cout(p_3_25[3]), .A(p_2_24[9]), .B(p_2_24[8]), .Cin(p_2_24[7]));
full_adder fa_3_24_4(.S(p_3_24[10]), .Cout(p_3_25[4]), .A(p_2_24[6]), .B(p_2_24[5]), .Cin(p_2_24[4]));
full_adder fa_3_24_5(.S(p_3_24[11]), .Cout(p_3_25[5]), .A(p_2_24[3]), .B(p_2_24[2]), .Cin(p_2_24[1]));
full_adder fa_3_25_0(.S(p_3_25[6]), .Cout(p_3_26[0]), .A(p_2_25[18]), .B(p_2_25[17]), .Cin(p_2_25[16]));
full_adder fa_3_25_1(.S(p_3_25[7]), .Cout(p_3_26[1]), .A(p_2_25[15]), .B(p_2_25[14]), .Cin(p_2_25[13]));
full_adder fa_3_25_2(.S(p_3_25[8]), .Cout(p_3_26[2]), .A(p_2_25[12]), .B(p_2_25[11]), .Cin(p_2_25[10]));
full_adder fa_3_25_3(.S(p_3_25[9]), .Cout(p_3_26[3]), .A(p_2_25[9]), .B(p_2_25[8]), .Cin(p_2_25[7]));
full_adder fa_3_25_4(.S(p_3_25[10]), .Cout(p_3_26[4]), .A(p_2_25[6]), .B(p_2_25[5]), .Cin(p_2_25[4]));
full_adder fa_3_25_5(.S(p_3_25[11]), .Cout(p_3_26[5]), .A(p_2_25[3]), .B(p_2_25[2]), .Cin(p_2_25[1]));
full_adder fa_3_26_0(.S(p_3_26[6]), .Cout(p_3_27[0]), .A(p_2_26[18]), .B(p_2_26[17]), .Cin(p_2_26[16]));
full_adder fa_3_26_1(.S(p_3_26[7]), .Cout(p_3_27[1]), .A(p_2_26[15]), .B(p_2_26[14]), .Cin(p_2_26[13]));
full_adder fa_3_26_2(.S(p_3_26[8]), .Cout(p_3_27[2]), .A(p_2_26[12]), .B(p_2_26[11]), .Cin(p_2_26[10]));
full_adder fa_3_26_3(.S(p_3_26[9]), .Cout(p_3_27[3]), .A(p_2_26[9]), .B(p_2_26[8]), .Cin(p_2_26[7]));
full_adder fa_3_26_4(.S(p_3_26[10]), .Cout(p_3_27[4]), .A(p_2_26[6]), .B(p_2_26[5]), .Cin(p_2_26[4]));
full_adder fa_3_26_5(.S(p_3_26[11]), .Cout(p_3_27[5]), .A(p_2_26[3]), .B(p_2_26[2]), .Cin(p_2_26[1]));
full_adder fa_3_27_0(.S(p_3_27[6]), .Cout(p_3_28[0]), .A(p_2_27[18]), .B(p_2_27[17]), .Cin(p_2_27[16]));
full_adder fa_3_27_1(.S(p_3_27[7]), .Cout(p_3_28[1]), .A(p_2_27[15]), .B(p_2_27[14]), .Cin(p_2_27[13]));
full_adder fa_3_27_2(.S(p_3_27[8]), .Cout(p_3_28[2]), .A(p_2_27[12]), .B(p_2_27[11]), .Cin(p_2_27[10]));
full_adder fa_3_27_3(.S(p_3_27[9]), .Cout(p_3_28[3]), .A(p_2_27[9]), .B(p_2_27[8]), .Cin(p_2_27[7]));
full_adder fa_3_27_4(.S(p_3_27[10]), .Cout(p_3_28[4]), .A(p_2_27[6]), .B(p_2_27[5]), .Cin(p_2_27[4]));
full_adder fa_3_27_5(.S(p_3_27[11]), .Cout(p_3_28[5]), .A(p_2_27[3]), .B(p_2_27[2]), .Cin(p_2_27[1]));
full_adder fa_3_28_0(.S(p_3_28[6]), .Cout(p_3_29[0]), .A(p_2_28[18]), .B(p_2_28[17]), .Cin(p_2_28[16]));
full_adder fa_3_28_1(.S(p_3_28[7]), .Cout(p_3_29[1]), .A(p_2_28[15]), .B(p_2_28[14]), .Cin(p_2_28[13]));
full_adder fa_3_28_2(.S(p_3_28[8]), .Cout(p_3_29[2]), .A(p_2_28[12]), .B(p_2_28[11]), .Cin(p_2_28[10]));
full_adder fa_3_28_3(.S(p_3_28[9]), .Cout(p_3_29[3]), .A(p_2_28[9]), .B(p_2_28[8]), .Cin(p_2_28[7]));
full_adder fa_3_28_4(.S(p_3_28[10]), .Cout(p_3_29[4]), .A(p_2_28[6]), .B(p_2_28[5]), .Cin(p_2_28[4]));
full_adder fa_3_28_5(.S(p_3_28[11]), .Cout(p_3_29[5]), .A(p_2_28[3]), .B(p_2_28[2]), .Cin(p_2_28[1]));
full_adder fa_3_29_0(.S(p_3_29[6]), .Cout(p_3_30[0]), .A(p_2_29[18]), .B(p_2_29[17]), .Cin(p_2_29[16]));
full_adder fa_3_29_1(.S(p_3_29[7]), .Cout(p_3_30[1]), .A(p_2_29[15]), .B(p_2_29[14]), .Cin(p_2_29[13]));
full_adder fa_3_29_2(.S(p_3_29[8]), .Cout(p_3_30[2]), .A(p_2_29[12]), .B(p_2_29[11]), .Cin(p_2_29[10]));
full_adder fa_3_29_3(.S(p_3_29[9]), .Cout(p_3_30[3]), .A(p_2_29[9]), .B(p_2_29[8]), .Cin(p_2_29[7]));
full_adder fa_3_29_4(.S(p_3_29[10]), .Cout(p_3_30[4]), .A(p_2_29[6]), .B(p_2_29[5]), .Cin(p_2_29[4]));
full_adder fa_3_29_5(.S(p_3_29[11]), .Cout(p_3_30[5]), .A(p_2_29[3]), .B(p_2_29[2]), .Cin(p_2_29[1]));
full_adder fa_3_30_0(.S(p_3_30[6]), .Cout(p_3_31[0]), .A(p_2_30[18]), .B(p_2_30[17]), .Cin(p_2_30[16]));
full_adder fa_3_30_1(.S(p_3_30[7]), .Cout(p_3_31[1]), .A(p_2_30[15]), .B(p_2_30[14]), .Cin(p_2_30[13]));
full_adder fa_3_30_2(.S(p_3_30[8]), .Cout(p_3_31[2]), .A(p_2_30[12]), .B(p_2_30[11]), .Cin(p_2_30[10]));
full_adder fa_3_30_3(.S(p_3_30[9]), .Cout(p_3_31[3]), .A(p_2_30[9]), .B(p_2_30[8]), .Cin(p_2_30[7]));
full_adder fa_3_30_4(.S(p_3_30[10]), .Cout(p_3_31[4]), .A(p_2_30[6]), .B(p_2_30[5]), .Cin(p_2_30[4]));
full_adder fa_3_30_5(.S(p_3_30[11]), .Cout(p_3_31[5]), .A(p_2_30[3]), .B(p_2_30[2]), .Cin(p_2_30[1]));
full_adder fa_3_31_0(.S(p_3_31[6]), .Cout(p_3_32[0]), .A(p_2_31[18]), .B(p_2_31[17]), .Cin(p_2_31[16]));
full_adder fa_3_31_1(.S(p_3_31[7]), .Cout(p_3_32[1]), .A(p_2_31[15]), .B(p_2_31[14]), .Cin(p_2_31[13]));
full_adder fa_3_31_2(.S(p_3_31[8]), .Cout(p_3_32[2]), .A(p_2_31[12]), .B(p_2_31[11]), .Cin(p_2_31[10]));
full_adder fa_3_31_3(.S(p_3_31[9]), .Cout(p_3_32[3]), .A(p_2_31[9]), .B(p_2_31[8]), .Cin(p_2_31[7]));
full_adder fa_3_31_4(.S(p_3_31[10]), .Cout(p_3_32[4]), .A(p_2_31[6]), .B(p_2_31[5]), .Cin(p_2_31[4]));
full_adder fa_3_31_5(.S(p_3_31[11]), .Cout(p_3_32[5]), .A(p_2_31[3]), .B(p_2_31[2]), .Cin(p_2_31[1]));
full_adder fa_3_32_0(.S(p_3_32[6]), .Cout(p_3_33[0]), .A(p_2_32[18]), .B(p_2_32[17]), .Cin(p_2_32[16]));
full_adder fa_3_32_1(.S(p_3_32[7]), .Cout(p_3_33[1]), .A(p_2_32[15]), .B(p_2_32[14]), .Cin(p_2_32[13]));
full_adder fa_3_32_2(.S(p_3_32[8]), .Cout(p_3_33[2]), .A(p_2_32[12]), .B(p_2_32[11]), .Cin(p_2_32[10]));
full_adder fa_3_32_3(.S(p_3_32[9]), .Cout(p_3_33[3]), .A(p_2_32[9]), .B(p_2_32[8]), .Cin(p_2_32[7]));
full_adder fa_3_32_4(.S(p_3_32[10]), .Cout(p_3_33[4]), .A(p_2_32[6]), .B(p_2_32[5]), .Cin(p_2_32[4]));
full_adder fa_3_32_5(.S(p_3_32[11]), .Cout(p_3_33[5]), .A(p_2_32[3]), .B(p_2_32[2]), .Cin(p_2_32[1]));
full_adder fa_3_33_0(.S(p_3_33[6]), .Cout(p_3_34[0]), .A(p_2_33[18]), .B(p_2_33[17]), .Cin(p_2_33[16]));
full_adder fa_3_33_1(.S(p_3_33[7]), .Cout(p_3_34[1]), .A(p_2_33[15]), .B(p_2_33[14]), .Cin(p_2_33[13]));
full_adder fa_3_33_2(.S(p_3_33[8]), .Cout(p_3_34[2]), .A(p_2_33[12]), .B(p_2_33[11]), .Cin(p_2_33[10]));
full_adder fa_3_33_3(.S(p_3_33[9]), .Cout(p_3_34[3]), .A(p_2_33[9]), .B(p_2_33[8]), .Cin(p_2_33[7]));
full_adder fa_3_33_4(.S(p_3_33[10]), .Cout(p_3_34[4]), .A(p_2_33[6]), .B(p_2_33[5]), .Cin(p_2_33[4]));
full_adder fa_3_33_5(.S(p_3_33[11]), .Cout(p_3_34[5]), .A(p_2_33[3]), .B(p_2_33[2]), .Cin(p_2_33[1]));
full_adder fa_3_34_0(.S(p_3_34[6]), .Cout(p_3_35[0]), .A(p_2_34[18]), .B(p_2_34[17]), .Cin(p_2_34[16]));
full_adder fa_3_34_1(.S(p_3_34[7]), .Cout(p_3_35[1]), .A(p_2_34[15]), .B(p_2_34[14]), .Cin(p_2_34[13]));
full_adder fa_3_34_2(.S(p_3_34[8]), .Cout(p_3_35[2]), .A(p_2_34[12]), .B(p_2_34[11]), .Cin(p_2_34[10]));
full_adder fa_3_34_3(.S(p_3_34[9]), .Cout(p_3_35[3]), .A(p_2_34[9]), .B(p_2_34[8]), .Cin(p_2_34[7]));
full_adder fa_3_34_4(.S(p_3_34[10]), .Cout(p_3_35[4]), .A(p_2_34[6]), .B(p_2_34[5]), .Cin(p_2_34[4]));
full_adder fa_3_34_5(.S(p_3_34[11]), .Cout(p_3_35[5]), .A(p_2_34[3]), .B(p_2_34[2]), .Cin(p_2_34[1]));
full_adder fa_3_35_0(.S(p_3_35[6]), .Cout(p_3_36[0]), .A(p_2_35[18]), .B(p_2_35[17]), .Cin(p_2_35[16]));
full_adder fa_3_35_1(.S(p_3_35[7]), .Cout(p_3_36[1]), .A(p_2_35[15]), .B(p_2_35[14]), .Cin(p_2_35[13]));
full_adder fa_3_35_2(.S(p_3_35[8]), .Cout(p_3_36[2]), .A(p_2_35[12]), .B(p_2_35[11]), .Cin(p_2_35[10]));
full_adder fa_3_35_3(.S(p_3_35[9]), .Cout(p_3_36[3]), .A(p_2_35[9]), .B(p_2_35[8]), .Cin(p_2_35[7]));
full_adder fa_3_35_4(.S(p_3_35[10]), .Cout(p_3_36[4]), .A(p_2_35[6]), .B(p_2_35[5]), .Cin(p_2_35[4]));
full_adder fa_3_35_5(.S(p_3_35[11]), .Cout(p_3_36[5]), .A(p_2_35[3]), .B(p_2_35[2]), .Cin(p_2_35[1]));
full_adder fa_3_36_0(.S(p_3_36[6]), .Cout(p_3_37[0]), .A(p_2_36[18]), .B(p_2_36[17]), .Cin(p_2_36[16]));
full_adder fa_3_36_1(.S(p_3_36[7]), .Cout(p_3_37[1]), .A(p_2_36[15]), .B(p_2_36[14]), .Cin(p_2_36[13]));
full_adder fa_3_36_2(.S(p_3_36[8]), .Cout(p_3_37[2]), .A(p_2_36[12]), .B(p_2_36[11]), .Cin(p_2_36[10]));
full_adder fa_3_36_3(.S(p_3_36[9]), .Cout(p_3_37[3]), .A(p_2_36[9]), .B(p_2_36[8]), .Cin(p_2_36[7]));
full_adder fa_3_36_4(.S(p_3_36[10]), .Cout(p_3_37[4]), .A(p_2_36[6]), .B(p_2_36[5]), .Cin(p_2_36[4]));
full_adder fa_3_36_5(.S(p_3_36[11]), .Cout(p_3_37[5]), .A(p_2_36[3]), .B(p_2_36[2]), .Cin(p_2_36[1]));
full_adder fa_3_37_0(.S(p_3_37[6]), .Cout(p_3_38[0]), .A(p_2_37[18]), .B(p_2_37[17]), .Cin(p_2_37[16]));
full_adder fa_3_37_1(.S(p_3_37[7]), .Cout(p_3_38[1]), .A(p_2_37[15]), .B(p_2_37[14]), .Cin(p_2_37[13]));
full_adder fa_3_37_2(.S(p_3_37[8]), .Cout(p_3_38[2]), .A(p_2_37[12]), .B(p_2_37[11]), .Cin(p_2_37[10]));
full_adder fa_3_37_3(.S(p_3_37[9]), .Cout(p_3_38[3]), .A(p_2_37[9]), .B(p_2_37[8]), .Cin(p_2_37[7]));
full_adder fa_3_37_4(.S(p_3_37[10]), .Cout(p_3_38[4]), .A(p_2_37[6]), .B(p_2_37[5]), .Cin(p_2_37[4]));
full_adder fa_3_37_5(.S(p_3_37[11]), .Cout(p_3_38[5]), .A(p_2_37[3]), .B(p_2_37[2]), .Cin(p_2_37[1]));
full_adder fa_3_38_0(.S(p_3_38[6]), .Cout(p_3_39[0]), .A(p_2_38[18]), .B(p_2_38[17]), .Cin(p_2_38[16]));
full_adder fa_3_38_1(.S(p_3_38[7]), .Cout(p_3_39[1]), .A(p_2_38[15]), .B(p_2_38[14]), .Cin(p_2_38[13]));
full_adder fa_3_38_2(.S(p_3_38[8]), .Cout(p_3_39[2]), .A(p_2_38[12]), .B(p_2_38[11]), .Cin(p_2_38[10]));
full_adder fa_3_38_3(.S(p_3_38[9]), .Cout(p_3_39[3]), .A(p_2_38[9]), .B(p_2_38[8]), .Cin(p_2_38[7]));
full_adder fa_3_38_4(.S(p_3_38[10]), .Cout(p_3_39[4]), .A(p_2_38[6]), .B(p_2_38[5]), .Cin(p_2_38[4]));
full_adder fa_3_38_5(.S(p_3_38[11]), .Cout(p_3_39[5]), .A(p_2_38[3]), .B(p_2_38[2]), .Cin(p_2_38[1]));
full_adder fa_3_39_0(.S(p_3_39[6]), .Cout(p_3_40[0]), .A(p_2_39[18]), .B(p_2_39[17]), .Cin(p_2_39[16]));
full_adder fa_3_39_1(.S(p_3_39[7]), .Cout(p_3_40[1]), .A(p_2_39[15]), .B(p_2_39[14]), .Cin(p_2_39[13]));
full_adder fa_3_39_2(.S(p_3_39[8]), .Cout(p_3_40[2]), .A(p_2_39[12]), .B(p_2_39[11]), .Cin(p_2_39[10]));
full_adder fa_3_39_3(.S(p_3_39[9]), .Cout(p_3_40[3]), .A(p_2_39[9]), .B(p_2_39[8]), .Cin(p_2_39[7]));
full_adder fa_3_39_4(.S(p_3_39[10]), .Cout(p_3_40[4]), .A(p_2_39[6]), .B(p_2_39[5]), .Cin(p_2_39[4]));
full_adder fa_3_39_5(.S(p_3_39[11]), .Cout(p_3_40[5]), .A(p_2_39[3]), .B(p_2_39[2]), .Cin(p_2_39[1]));
full_adder fa_3_40_0(.S(p_3_40[6]), .Cout(p_3_41[0]), .A(p_2_40[18]), .B(p_2_40[17]), .Cin(p_2_40[16]));
full_adder fa_3_40_1(.S(p_3_40[7]), .Cout(p_3_41[1]), .A(p_2_40[15]), .B(p_2_40[14]), .Cin(p_2_40[13]));
full_adder fa_3_40_2(.S(p_3_40[8]), .Cout(p_3_41[2]), .A(p_2_40[12]), .B(p_2_40[11]), .Cin(p_2_40[10]));
full_adder fa_3_40_3(.S(p_3_40[9]), .Cout(p_3_41[3]), .A(p_2_40[9]), .B(p_2_40[8]), .Cin(p_2_40[7]));
full_adder fa_3_40_4(.S(p_3_40[10]), .Cout(p_3_41[4]), .A(p_2_40[6]), .B(p_2_40[5]), .Cin(p_2_40[4]));
full_adder fa_3_40_5(.S(p_3_40[11]), .Cout(p_3_41[5]), .A(p_2_40[3]), .B(p_2_40[2]), .Cin(p_2_40[1]));
full_adder fa_3_41_0(.S(p_3_41[6]), .Cout(p_3_42[0]), .A(p_2_41[18]), .B(p_2_41[17]), .Cin(p_2_41[16]));
full_adder fa_3_41_1(.S(p_3_41[7]), .Cout(p_3_42[1]), .A(p_2_41[15]), .B(p_2_41[14]), .Cin(p_2_41[13]));
full_adder fa_3_41_2(.S(p_3_41[8]), .Cout(p_3_42[2]), .A(p_2_41[12]), .B(p_2_41[11]), .Cin(p_2_41[10]));
full_adder fa_3_41_3(.S(p_3_41[9]), .Cout(p_3_42[3]), .A(p_2_41[9]), .B(p_2_41[8]), .Cin(p_2_41[7]));
full_adder fa_3_41_4(.S(p_3_41[10]), .Cout(p_3_42[4]), .A(p_2_41[6]), .B(p_2_41[5]), .Cin(p_2_41[4]));
full_adder fa_3_41_5(.S(p_3_41[11]), .Cout(p_3_42[5]), .A(p_2_41[3]), .B(p_2_41[2]), .Cin(p_2_41[1]));
full_adder fa_3_42_0(.S(p_3_42[6]), .Cout(p_3_43[0]), .A(p_2_42[18]), .B(p_2_42[17]), .Cin(p_2_42[16]));
full_adder fa_3_42_1(.S(p_3_42[7]), .Cout(p_3_43[1]), .A(p_2_42[15]), .B(p_2_42[14]), .Cin(p_2_42[13]));
full_adder fa_3_42_2(.S(p_3_42[8]), .Cout(p_3_43[2]), .A(p_2_42[12]), .B(p_2_42[11]), .Cin(p_2_42[10]));
full_adder fa_3_42_3(.S(p_3_42[9]), .Cout(p_3_43[3]), .A(p_2_42[9]), .B(p_2_42[8]), .Cin(p_2_42[7]));
full_adder fa_3_42_4(.S(p_3_42[10]), .Cout(p_3_43[4]), .A(p_2_42[6]), .B(p_2_42[5]), .Cin(p_2_42[4]));
full_adder fa_3_42_5(.S(p_3_42[11]), .Cout(p_3_43[5]), .A(p_2_42[3]), .B(p_2_42[2]), .Cin(p_2_42[1]));
full_adder fa_3_43_0(.S(p_3_43[6]), .Cout(p_3_44[0]), .A(p_2_43[18]), .B(p_2_43[17]), .Cin(p_2_43[16]));
full_adder fa_3_43_1(.S(p_3_43[7]), .Cout(p_3_44[1]), .A(p_2_43[15]), .B(p_2_43[14]), .Cin(p_2_43[13]));
full_adder fa_3_43_2(.S(p_3_43[8]), .Cout(p_3_44[2]), .A(p_2_43[12]), .B(p_2_43[11]), .Cin(p_2_43[10]));
full_adder fa_3_43_3(.S(p_3_43[9]), .Cout(p_3_44[3]), .A(p_2_43[9]), .B(p_2_43[8]), .Cin(p_2_43[7]));
full_adder fa_3_43_4(.S(p_3_43[10]), .Cout(p_3_44[4]), .A(p_2_43[6]), .B(p_2_43[5]), .Cin(p_2_43[4]));
full_adder fa_3_43_5(.S(p_3_43[11]), .Cout(p_3_44[5]), .A(p_2_43[3]), .B(p_2_43[2]), .Cin(p_2_43[1]));
full_adder fa_3_44_0(.S(p_3_44[6]), .Cout(p_3_45[0]), .A(p_2_44[18]), .B(p_2_44[17]), .Cin(p_2_44[16]));
full_adder fa_3_44_1(.S(p_3_44[7]), .Cout(p_3_45[1]), .A(p_2_44[15]), .B(p_2_44[14]), .Cin(p_2_44[13]));
full_adder fa_3_44_2(.S(p_3_44[8]), .Cout(p_3_45[2]), .A(p_2_44[12]), .B(p_2_44[11]), .Cin(p_2_44[10]));
full_adder fa_3_44_3(.S(p_3_44[9]), .Cout(p_3_45[3]), .A(p_2_44[9]), .B(p_2_44[8]), .Cin(p_2_44[7]));
full_adder fa_3_44_4(.S(p_3_44[10]), .Cout(p_3_45[4]), .A(p_2_44[6]), .B(p_2_44[5]), .Cin(p_2_44[4]));
full_adder fa_3_44_5(.S(p_3_44[11]), .Cout(p_3_45[5]), .A(p_2_44[3]), .B(p_2_44[2]), .Cin(p_2_44[1]));
full_adder fa_3_45_0(.S(p_3_45[6]), .Cout(p_3_46[0]), .A(p_2_45[18]), .B(p_2_45[17]), .Cin(p_2_45[16]));
full_adder fa_3_45_1(.S(p_3_45[7]), .Cout(p_3_46[1]), .A(p_2_45[15]), .B(p_2_45[14]), .Cin(p_2_45[13]));
full_adder fa_3_45_2(.S(p_3_45[8]), .Cout(p_3_46[2]), .A(p_2_45[12]), .B(p_2_45[11]), .Cin(p_2_45[10]));
full_adder fa_3_45_3(.S(p_3_45[9]), .Cout(p_3_46[3]), .A(p_2_45[9]), .B(p_2_45[8]), .Cin(p_2_45[7]));
full_adder fa_3_45_4(.S(p_3_45[10]), .Cout(p_3_46[4]), .A(p_2_45[6]), .B(p_2_45[5]), .Cin(p_2_45[4]));
full_adder fa_3_45_5(.S(p_3_45[11]), .Cout(p_3_46[5]), .A(p_2_45[3]), .B(p_2_45[2]), .Cin(p_2_45[1]));
full_adder fa_3_46_0(.S(p_3_46[6]), .Cout(p_3_47[0]), .A(p_2_46[16]), .B(p_2_46[15]), .Cin(p_2_46[14]));
full_adder fa_3_46_1(.S(p_3_46[7]), .Cout(p_3_47[1]), .A(p_2_46[13]), .B(p_2_46[12]), .Cin(p_2_46[11]));
full_adder fa_3_46_2(.S(p_3_46[8]), .Cout(p_3_47[2]), .A(p_2_46[10]), .B(p_2_46[9]), .Cin(p_2_46[8]));
full_adder fa_3_46_3(.S(p_3_46[9]), .Cout(p_3_47[3]), .A(p_2_46[7]), .B(p_2_46[6]), .Cin(p_2_46[5]));
full_adder fa_3_46_4(.S(p_3_46[10]), .Cout(p_3_47[4]), .A(p_2_46[4]), .B(p_2_46[3]), .Cin(p_2_46[2]));
full_adder fa_3_47_0(.S(p_3_47[5]), .Cout(p_3_48[0]), .A(p_2_47[15]), .B(p_2_47[14]), .Cin(p_2_47[13]));
full_adder fa_3_47_1(.S(p_3_47[6]), .Cout(p_3_48[1]), .A(p_2_47[12]), .B(p_2_47[11]), .Cin(p_2_47[10]));
full_adder fa_3_47_2(.S(p_3_47[7]), .Cout(p_3_48[2]), .A(p_2_47[9]), .B(p_2_47[8]), .Cin(p_2_47[7]));
full_adder fa_3_47_3(.S(p_3_47[8]), .Cout(p_3_48[3]), .A(p_2_47[6]), .B(p_2_47[5]), .Cin(p_2_47[4]));
full_adder fa_3_48_0(.S(p_3_48[4]), .Cout(p_3_49[0]), .A(p_2_48[14]), .B(p_2_48[13]), .Cin(p_2_48[12]));
full_adder fa_3_48_1(.S(p_3_48[5]), .Cout(p_3_49[1]), .A(p_2_48[11]), .B(p_2_48[10]), .Cin(p_2_48[9]));
full_adder fa_3_48_2(.S(p_3_48[6]), .Cout(p_3_49[2]), .A(p_2_48[8]), .B(p_2_48[7]), .Cin(p_2_48[6]));
full_adder fa_3_49_0(.S(p_3_49[3]), .Cout(p_3_50[0]), .A(p_2_49[13]), .B(p_2_49[12]), .Cin(p_2_49[11]));
full_adder fa_3_49_1(.S(p_3_49[4]), .Cout(p_3_50[1]), .A(p_2_49[10]), .B(p_2_49[9]), .Cin(p_2_49[8]));
full_adder fa_3_50_0(.S(p_3_50[2]), .Cout(p_3_51[0]), .A(p_2_50[12]), .B(p_2_50[11]), .Cin(p_2_50[10]));

// Stage 4 non-added partial products
assign p_4_0[0:0] = p_3_0[0:0];
assign p_4_1[1:0] = p_3_1[1:0];
assign p_4_2[2:0] = p_3_2[2:0];
assign p_4_3[3:0] = p_3_3[3:0];
assign p_4_4[4:0] = p_3_4[4:0];
assign p_4_5[5:0] = p_3_5[5:0];
assign p_4_6[6:0] = p_3_6[6:0];
assign p_4_7[7:0] = p_3_7[7:0];
assign p_4_8[8:0] = p_3_8[8:0];
assign p_4_9[8:1] = p_3_9[7:0];
assign p_4_10[8:3] = p_3_10[5:0];
assign p_4_11[8:5] = p_3_11[3:0];
assign p_4_12[8:7] = p_3_12[1:0];
assign p_4_13[8:8] = p_3_13[0:0];
assign p_4_14[8:8] = p_3_14[0:0];
assign p_4_15[8:8] = p_3_15[0:0];
assign p_4_16[8:8] = p_3_16[0:0];
assign p_4_17[8:8] = p_3_17[0:0];
assign p_4_18[8:8] = p_3_18[0:0];
assign p_4_19[8:8] = p_3_19[0:0];
assign p_4_20[8:8] = p_3_20[0:0];
assign p_4_21[8:8] = p_3_21[0:0];
assign p_4_22[8:8] = p_3_22[0:0];
assign p_4_23[8:8] = p_3_23[0:0];
assign p_4_24[8:8] = p_3_24[0:0];
assign p_4_25[8:8] = p_3_25[0:0];
assign p_4_26[8:8] = p_3_26[0:0];
assign p_4_27[8:8] = p_3_27[0:0];
assign p_4_28[8:8] = p_3_28[0:0];
assign p_4_29[8:8] = p_3_29[0:0];
assign p_4_30[8:8] = p_3_30[0:0];
assign p_4_31[8:8] = p_3_31[0:0];
assign p_4_32[8:8] = p_3_32[0:0];
assign p_4_33[8:8] = p_3_33[0:0];
assign p_4_34[8:8] = p_3_34[0:0];
assign p_4_35[8:8] = p_3_35[0:0];
assign p_4_36[8:8] = p_3_36[0:0];
assign p_4_37[8:8] = p_3_37[0:0];
assign p_4_38[8:8] = p_3_38[0:0];
assign p_4_39[8:8] = p_3_39[0:0];
assign p_4_40[8:8] = p_3_40[0:0];
assign p_4_41[8:8] = p_3_41[0:0];
assign p_4_42[8:8] = p_3_42[0:0];
assign p_4_43[8:8] = p_3_43[0:0];
assign p_4_44[8:8] = p_3_44[0:0];
assign p_4_45[8:8] = p_3_45[0:0];
assign p_4_46[8:8] = p_3_46[0:0];
assign p_4_47[8:8] = p_3_47[0:0];
assign p_4_48[8:8] = p_3_48[0:0];
assign p_4_49[8:8] = p_3_49[0:0];
assign p_4_50[8:8] = p_3_50[0:0];
assign p_4_51[8:8] = p_3_51[0:0];
assign p_4_52[8:7] = p_3_52[1:0];
assign p_4_53[8:5] = p_3_53[3:0];
assign p_4_54[8:3] = p_3_54[5:0];
assign p_4_55[8:1] = p_3_55[7:0];
assign p_4_56[6:0] = p_3_56[6:0];
assign p_4_57[5:0] = p_3_57[5:0];
assign p_4_58[4:0] = p_3_58[4:0];
assign p_4_59[3:0] = p_3_59[3:0];
assign p_4_60[2:0] = p_3_60[2:0];
assign p_4_61[1:0] = p_3_61[1:0];
assign p_4_62[0:0] = p_3_62[0:0];
// Stage 4 adders
half_adder ha_4_9(.S(p_4_9[0]), .Cout(p_4_10[0]), .A(p_3_9[9]), .B(p_3_9[8]));
full_adder fa_4_10_0(.S(p_4_10[1]), .Cout(p_4_11[0]), .A(p_3_10[10]), .B(p_3_10[9]), .Cin(p_3_10[8]));
half_adder ha_4_10(.S(p_4_10[2]), .Cout(p_4_11[1]), .A(p_3_10[7]), .B(p_3_10[6]));
full_adder fa_4_11_0(.S(p_4_11[2]), .Cout(p_4_12[0]), .A(p_3_11[11]), .B(p_3_11[10]), .Cin(p_3_11[9]));
full_adder fa_4_11_1(.S(p_4_11[3]), .Cout(p_4_12[1]), .A(p_3_11[8]), .B(p_3_11[7]), .Cin(p_3_11[6]));
half_adder ha_4_11(.S(p_4_11[4]), .Cout(p_4_12[2]), .A(p_3_11[5]), .B(p_3_11[4]));
full_adder fa_4_12_0(.S(p_4_12[3]), .Cout(p_4_13[0]), .A(p_3_12[12]), .B(p_3_12[11]), .Cin(p_3_12[10]));
full_adder fa_4_12_1(.S(p_4_12[4]), .Cout(p_4_13[1]), .A(p_3_12[9]), .B(p_3_12[8]), .Cin(p_3_12[7]));
full_adder fa_4_12_2(.S(p_4_12[5]), .Cout(p_4_13[2]), .A(p_3_12[6]), .B(p_3_12[5]), .Cin(p_3_12[4]));
half_adder ha_4_12(.S(p_4_12[6]), .Cout(p_4_13[3]), .A(p_3_12[3]), .B(p_3_12[2]));
full_adder fa_4_13_0(.S(p_4_13[4]), .Cout(p_4_14[0]), .A(p_3_13[12]), .B(p_3_13[11]), .Cin(p_3_13[10]));
full_adder fa_4_13_1(.S(p_4_13[5]), .Cout(p_4_14[1]), .A(p_3_13[9]), .B(p_3_13[8]), .Cin(p_3_13[7]));
full_adder fa_4_13_2(.S(p_4_13[6]), .Cout(p_4_14[2]), .A(p_3_13[6]), .B(p_3_13[5]), .Cin(p_3_13[4]));
full_adder fa_4_13_3(.S(p_4_13[7]), .Cout(p_4_14[3]), .A(p_3_13[3]), .B(p_3_13[2]), .Cin(p_3_13[1]));
full_adder fa_4_14_0(.S(p_4_14[4]), .Cout(p_4_15[0]), .A(p_3_14[12]), .B(p_3_14[11]), .Cin(p_3_14[10]));
full_adder fa_4_14_1(.S(p_4_14[5]), .Cout(p_4_15[1]), .A(p_3_14[9]), .B(p_3_14[8]), .Cin(p_3_14[7]));
full_adder fa_4_14_2(.S(p_4_14[6]), .Cout(p_4_15[2]), .A(p_3_14[6]), .B(p_3_14[5]), .Cin(p_3_14[4]));
full_adder fa_4_14_3(.S(p_4_14[7]), .Cout(p_4_15[3]), .A(p_3_14[3]), .B(p_3_14[2]), .Cin(p_3_14[1]));
full_adder fa_4_15_0(.S(p_4_15[4]), .Cout(p_4_16[0]), .A(p_3_15[12]), .B(p_3_15[11]), .Cin(p_3_15[10]));
full_adder fa_4_15_1(.S(p_4_15[5]), .Cout(p_4_16[1]), .A(p_3_15[9]), .B(p_3_15[8]), .Cin(p_3_15[7]));
full_adder fa_4_15_2(.S(p_4_15[6]), .Cout(p_4_16[2]), .A(p_3_15[6]), .B(p_3_15[5]), .Cin(p_3_15[4]));
full_adder fa_4_15_3(.S(p_4_15[7]), .Cout(p_4_16[3]), .A(p_3_15[3]), .B(p_3_15[2]), .Cin(p_3_15[1]));
full_adder fa_4_16_0(.S(p_4_16[4]), .Cout(p_4_17[0]), .A(p_3_16[12]), .B(p_3_16[11]), .Cin(p_3_16[10]));
full_adder fa_4_16_1(.S(p_4_16[5]), .Cout(p_4_17[1]), .A(p_3_16[9]), .B(p_3_16[8]), .Cin(p_3_16[7]));
full_adder fa_4_16_2(.S(p_4_16[6]), .Cout(p_4_17[2]), .A(p_3_16[6]), .B(p_3_16[5]), .Cin(p_3_16[4]));
full_adder fa_4_16_3(.S(p_4_16[7]), .Cout(p_4_17[3]), .A(p_3_16[3]), .B(p_3_16[2]), .Cin(p_3_16[1]));
full_adder fa_4_17_0(.S(p_4_17[4]), .Cout(p_4_18[0]), .A(p_3_17[12]), .B(p_3_17[11]), .Cin(p_3_17[10]));
full_adder fa_4_17_1(.S(p_4_17[5]), .Cout(p_4_18[1]), .A(p_3_17[9]), .B(p_3_17[8]), .Cin(p_3_17[7]));
full_adder fa_4_17_2(.S(p_4_17[6]), .Cout(p_4_18[2]), .A(p_3_17[6]), .B(p_3_17[5]), .Cin(p_3_17[4]));
full_adder fa_4_17_3(.S(p_4_17[7]), .Cout(p_4_18[3]), .A(p_3_17[3]), .B(p_3_17[2]), .Cin(p_3_17[1]));
full_adder fa_4_18_0(.S(p_4_18[4]), .Cout(p_4_19[0]), .A(p_3_18[12]), .B(p_3_18[11]), .Cin(p_3_18[10]));
full_adder fa_4_18_1(.S(p_4_18[5]), .Cout(p_4_19[1]), .A(p_3_18[9]), .B(p_3_18[8]), .Cin(p_3_18[7]));
full_adder fa_4_18_2(.S(p_4_18[6]), .Cout(p_4_19[2]), .A(p_3_18[6]), .B(p_3_18[5]), .Cin(p_3_18[4]));
full_adder fa_4_18_3(.S(p_4_18[7]), .Cout(p_4_19[3]), .A(p_3_18[3]), .B(p_3_18[2]), .Cin(p_3_18[1]));
full_adder fa_4_19_0(.S(p_4_19[4]), .Cout(p_4_20[0]), .A(p_3_19[12]), .B(p_3_19[11]), .Cin(p_3_19[10]));
full_adder fa_4_19_1(.S(p_4_19[5]), .Cout(p_4_20[1]), .A(p_3_19[9]), .B(p_3_19[8]), .Cin(p_3_19[7]));
full_adder fa_4_19_2(.S(p_4_19[6]), .Cout(p_4_20[2]), .A(p_3_19[6]), .B(p_3_19[5]), .Cin(p_3_19[4]));
full_adder fa_4_19_3(.S(p_4_19[7]), .Cout(p_4_20[3]), .A(p_3_19[3]), .B(p_3_19[2]), .Cin(p_3_19[1]));
full_adder fa_4_20_0(.S(p_4_20[4]), .Cout(p_4_21[0]), .A(p_3_20[12]), .B(p_3_20[11]), .Cin(p_3_20[10]));
full_adder fa_4_20_1(.S(p_4_20[5]), .Cout(p_4_21[1]), .A(p_3_20[9]), .B(p_3_20[8]), .Cin(p_3_20[7]));
full_adder fa_4_20_2(.S(p_4_20[6]), .Cout(p_4_21[2]), .A(p_3_20[6]), .B(p_3_20[5]), .Cin(p_3_20[4]));
full_adder fa_4_20_3(.S(p_4_20[7]), .Cout(p_4_21[3]), .A(p_3_20[3]), .B(p_3_20[2]), .Cin(p_3_20[1]));
full_adder fa_4_21_0(.S(p_4_21[4]), .Cout(p_4_22[0]), .A(p_3_21[12]), .B(p_3_21[11]), .Cin(p_3_21[10]));
full_adder fa_4_21_1(.S(p_4_21[5]), .Cout(p_4_22[1]), .A(p_3_21[9]), .B(p_3_21[8]), .Cin(p_3_21[7]));
full_adder fa_4_21_2(.S(p_4_21[6]), .Cout(p_4_22[2]), .A(p_3_21[6]), .B(p_3_21[5]), .Cin(p_3_21[4]));
full_adder fa_4_21_3(.S(p_4_21[7]), .Cout(p_4_22[3]), .A(p_3_21[3]), .B(p_3_21[2]), .Cin(p_3_21[1]));
full_adder fa_4_22_0(.S(p_4_22[4]), .Cout(p_4_23[0]), .A(p_3_22[12]), .B(p_3_22[11]), .Cin(p_3_22[10]));
full_adder fa_4_22_1(.S(p_4_22[5]), .Cout(p_4_23[1]), .A(p_3_22[9]), .B(p_3_22[8]), .Cin(p_3_22[7]));
full_adder fa_4_22_2(.S(p_4_22[6]), .Cout(p_4_23[2]), .A(p_3_22[6]), .B(p_3_22[5]), .Cin(p_3_22[4]));
full_adder fa_4_22_3(.S(p_4_22[7]), .Cout(p_4_23[3]), .A(p_3_22[3]), .B(p_3_22[2]), .Cin(p_3_22[1]));
full_adder fa_4_23_0(.S(p_4_23[4]), .Cout(p_4_24[0]), .A(p_3_23[12]), .B(p_3_23[11]), .Cin(p_3_23[10]));
full_adder fa_4_23_1(.S(p_4_23[5]), .Cout(p_4_24[1]), .A(p_3_23[9]), .B(p_3_23[8]), .Cin(p_3_23[7]));
full_adder fa_4_23_2(.S(p_4_23[6]), .Cout(p_4_24[2]), .A(p_3_23[6]), .B(p_3_23[5]), .Cin(p_3_23[4]));
full_adder fa_4_23_3(.S(p_4_23[7]), .Cout(p_4_24[3]), .A(p_3_23[3]), .B(p_3_23[2]), .Cin(p_3_23[1]));
full_adder fa_4_24_0(.S(p_4_24[4]), .Cout(p_4_25[0]), .A(p_3_24[12]), .B(p_3_24[11]), .Cin(p_3_24[10]));
full_adder fa_4_24_1(.S(p_4_24[5]), .Cout(p_4_25[1]), .A(p_3_24[9]), .B(p_3_24[8]), .Cin(p_3_24[7]));
full_adder fa_4_24_2(.S(p_4_24[6]), .Cout(p_4_25[2]), .A(p_3_24[6]), .B(p_3_24[5]), .Cin(p_3_24[4]));
full_adder fa_4_24_3(.S(p_4_24[7]), .Cout(p_4_25[3]), .A(p_3_24[3]), .B(p_3_24[2]), .Cin(p_3_24[1]));
full_adder fa_4_25_0(.S(p_4_25[4]), .Cout(p_4_26[0]), .A(p_3_25[12]), .B(p_3_25[11]), .Cin(p_3_25[10]));
full_adder fa_4_25_1(.S(p_4_25[5]), .Cout(p_4_26[1]), .A(p_3_25[9]), .B(p_3_25[8]), .Cin(p_3_25[7]));
full_adder fa_4_25_2(.S(p_4_25[6]), .Cout(p_4_26[2]), .A(p_3_25[6]), .B(p_3_25[5]), .Cin(p_3_25[4]));
full_adder fa_4_25_3(.S(p_4_25[7]), .Cout(p_4_26[3]), .A(p_3_25[3]), .B(p_3_25[2]), .Cin(p_3_25[1]));
full_adder fa_4_26_0(.S(p_4_26[4]), .Cout(p_4_27[0]), .A(p_3_26[12]), .B(p_3_26[11]), .Cin(p_3_26[10]));
full_adder fa_4_26_1(.S(p_4_26[5]), .Cout(p_4_27[1]), .A(p_3_26[9]), .B(p_3_26[8]), .Cin(p_3_26[7]));
full_adder fa_4_26_2(.S(p_4_26[6]), .Cout(p_4_27[2]), .A(p_3_26[6]), .B(p_3_26[5]), .Cin(p_3_26[4]));
full_adder fa_4_26_3(.S(p_4_26[7]), .Cout(p_4_27[3]), .A(p_3_26[3]), .B(p_3_26[2]), .Cin(p_3_26[1]));
full_adder fa_4_27_0(.S(p_4_27[4]), .Cout(p_4_28[0]), .A(p_3_27[12]), .B(p_3_27[11]), .Cin(p_3_27[10]));
full_adder fa_4_27_1(.S(p_4_27[5]), .Cout(p_4_28[1]), .A(p_3_27[9]), .B(p_3_27[8]), .Cin(p_3_27[7]));
full_adder fa_4_27_2(.S(p_4_27[6]), .Cout(p_4_28[2]), .A(p_3_27[6]), .B(p_3_27[5]), .Cin(p_3_27[4]));
full_adder fa_4_27_3(.S(p_4_27[7]), .Cout(p_4_28[3]), .A(p_3_27[3]), .B(p_3_27[2]), .Cin(p_3_27[1]));
full_adder fa_4_28_0(.S(p_4_28[4]), .Cout(p_4_29[0]), .A(p_3_28[12]), .B(p_3_28[11]), .Cin(p_3_28[10]));
full_adder fa_4_28_1(.S(p_4_28[5]), .Cout(p_4_29[1]), .A(p_3_28[9]), .B(p_3_28[8]), .Cin(p_3_28[7]));
full_adder fa_4_28_2(.S(p_4_28[6]), .Cout(p_4_29[2]), .A(p_3_28[6]), .B(p_3_28[5]), .Cin(p_3_28[4]));
full_adder fa_4_28_3(.S(p_4_28[7]), .Cout(p_4_29[3]), .A(p_3_28[3]), .B(p_3_28[2]), .Cin(p_3_28[1]));
full_adder fa_4_29_0(.S(p_4_29[4]), .Cout(p_4_30[0]), .A(p_3_29[12]), .B(p_3_29[11]), .Cin(p_3_29[10]));
full_adder fa_4_29_1(.S(p_4_29[5]), .Cout(p_4_30[1]), .A(p_3_29[9]), .B(p_3_29[8]), .Cin(p_3_29[7]));
full_adder fa_4_29_2(.S(p_4_29[6]), .Cout(p_4_30[2]), .A(p_3_29[6]), .B(p_3_29[5]), .Cin(p_3_29[4]));
full_adder fa_4_29_3(.S(p_4_29[7]), .Cout(p_4_30[3]), .A(p_3_29[3]), .B(p_3_29[2]), .Cin(p_3_29[1]));
full_adder fa_4_30_0(.S(p_4_30[4]), .Cout(p_4_31[0]), .A(p_3_30[12]), .B(p_3_30[11]), .Cin(p_3_30[10]));
full_adder fa_4_30_1(.S(p_4_30[5]), .Cout(p_4_31[1]), .A(p_3_30[9]), .B(p_3_30[8]), .Cin(p_3_30[7]));
full_adder fa_4_30_2(.S(p_4_30[6]), .Cout(p_4_31[2]), .A(p_3_30[6]), .B(p_3_30[5]), .Cin(p_3_30[4]));
full_adder fa_4_30_3(.S(p_4_30[7]), .Cout(p_4_31[3]), .A(p_3_30[3]), .B(p_3_30[2]), .Cin(p_3_30[1]));
full_adder fa_4_31_0(.S(p_4_31[4]), .Cout(p_4_32[0]), .A(p_3_31[12]), .B(p_3_31[11]), .Cin(p_3_31[10]));
full_adder fa_4_31_1(.S(p_4_31[5]), .Cout(p_4_32[1]), .A(p_3_31[9]), .B(p_3_31[8]), .Cin(p_3_31[7]));
full_adder fa_4_31_2(.S(p_4_31[6]), .Cout(p_4_32[2]), .A(p_3_31[6]), .B(p_3_31[5]), .Cin(p_3_31[4]));
full_adder fa_4_31_3(.S(p_4_31[7]), .Cout(p_4_32[3]), .A(p_3_31[3]), .B(p_3_31[2]), .Cin(p_3_31[1]));
full_adder fa_4_32_0(.S(p_4_32[4]), .Cout(p_4_33[0]), .A(p_3_32[12]), .B(p_3_32[11]), .Cin(p_3_32[10]));
full_adder fa_4_32_1(.S(p_4_32[5]), .Cout(p_4_33[1]), .A(p_3_32[9]), .B(p_3_32[8]), .Cin(p_3_32[7]));
full_adder fa_4_32_2(.S(p_4_32[6]), .Cout(p_4_33[2]), .A(p_3_32[6]), .B(p_3_32[5]), .Cin(p_3_32[4]));
full_adder fa_4_32_3(.S(p_4_32[7]), .Cout(p_4_33[3]), .A(p_3_32[3]), .B(p_3_32[2]), .Cin(p_3_32[1]));
full_adder fa_4_33_0(.S(p_4_33[4]), .Cout(p_4_34[0]), .A(p_3_33[12]), .B(p_3_33[11]), .Cin(p_3_33[10]));
full_adder fa_4_33_1(.S(p_4_33[5]), .Cout(p_4_34[1]), .A(p_3_33[9]), .B(p_3_33[8]), .Cin(p_3_33[7]));
full_adder fa_4_33_2(.S(p_4_33[6]), .Cout(p_4_34[2]), .A(p_3_33[6]), .B(p_3_33[5]), .Cin(p_3_33[4]));
full_adder fa_4_33_3(.S(p_4_33[7]), .Cout(p_4_34[3]), .A(p_3_33[3]), .B(p_3_33[2]), .Cin(p_3_33[1]));
full_adder fa_4_34_0(.S(p_4_34[4]), .Cout(p_4_35[0]), .A(p_3_34[12]), .B(p_3_34[11]), .Cin(p_3_34[10]));
full_adder fa_4_34_1(.S(p_4_34[5]), .Cout(p_4_35[1]), .A(p_3_34[9]), .B(p_3_34[8]), .Cin(p_3_34[7]));
full_adder fa_4_34_2(.S(p_4_34[6]), .Cout(p_4_35[2]), .A(p_3_34[6]), .B(p_3_34[5]), .Cin(p_3_34[4]));
full_adder fa_4_34_3(.S(p_4_34[7]), .Cout(p_4_35[3]), .A(p_3_34[3]), .B(p_3_34[2]), .Cin(p_3_34[1]));
full_adder fa_4_35_0(.S(p_4_35[4]), .Cout(p_4_36[0]), .A(p_3_35[12]), .B(p_3_35[11]), .Cin(p_3_35[10]));
full_adder fa_4_35_1(.S(p_4_35[5]), .Cout(p_4_36[1]), .A(p_3_35[9]), .B(p_3_35[8]), .Cin(p_3_35[7]));
full_adder fa_4_35_2(.S(p_4_35[6]), .Cout(p_4_36[2]), .A(p_3_35[6]), .B(p_3_35[5]), .Cin(p_3_35[4]));
full_adder fa_4_35_3(.S(p_4_35[7]), .Cout(p_4_36[3]), .A(p_3_35[3]), .B(p_3_35[2]), .Cin(p_3_35[1]));
full_adder fa_4_36_0(.S(p_4_36[4]), .Cout(p_4_37[0]), .A(p_3_36[12]), .B(p_3_36[11]), .Cin(p_3_36[10]));
full_adder fa_4_36_1(.S(p_4_36[5]), .Cout(p_4_37[1]), .A(p_3_36[9]), .B(p_3_36[8]), .Cin(p_3_36[7]));
full_adder fa_4_36_2(.S(p_4_36[6]), .Cout(p_4_37[2]), .A(p_3_36[6]), .B(p_3_36[5]), .Cin(p_3_36[4]));
full_adder fa_4_36_3(.S(p_4_36[7]), .Cout(p_4_37[3]), .A(p_3_36[3]), .B(p_3_36[2]), .Cin(p_3_36[1]));
full_adder fa_4_37_0(.S(p_4_37[4]), .Cout(p_4_38[0]), .A(p_3_37[12]), .B(p_3_37[11]), .Cin(p_3_37[10]));
full_adder fa_4_37_1(.S(p_4_37[5]), .Cout(p_4_38[1]), .A(p_3_37[9]), .B(p_3_37[8]), .Cin(p_3_37[7]));
full_adder fa_4_37_2(.S(p_4_37[6]), .Cout(p_4_38[2]), .A(p_3_37[6]), .B(p_3_37[5]), .Cin(p_3_37[4]));
full_adder fa_4_37_3(.S(p_4_37[7]), .Cout(p_4_38[3]), .A(p_3_37[3]), .B(p_3_37[2]), .Cin(p_3_37[1]));
full_adder fa_4_38_0(.S(p_4_38[4]), .Cout(p_4_39[0]), .A(p_3_38[12]), .B(p_3_38[11]), .Cin(p_3_38[10]));
full_adder fa_4_38_1(.S(p_4_38[5]), .Cout(p_4_39[1]), .A(p_3_38[9]), .B(p_3_38[8]), .Cin(p_3_38[7]));
full_adder fa_4_38_2(.S(p_4_38[6]), .Cout(p_4_39[2]), .A(p_3_38[6]), .B(p_3_38[5]), .Cin(p_3_38[4]));
full_adder fa_4_38_3(.S(p_4_38[7]), .Cout(p_4_39[3]), .A(p_3_38[3]), .B(p_3_38[2]), .Cin(p_3_38[1]));
full_adder fa_4_39_0(.S(p_4_39[4]), .Cout(p_4_40[0]), .A(p_3_39[12]), .B(p_3_39[11]), .Cin(p_3_39[10]));
full_adder fa_4_39_1(.S(p_4_39[5]), .Cout(p_4_40[1]), .A(p_3_39[9]), .B(p_3_39[8]), .Cin(p_3_39[7]));
full_adder fa_4_39_2(.S(p_4_39[6]), .Cout(p_4_40[2]), .A(p_3_39[6]), .B(p_3_39[5]), .Cin(p_3_39[4]));
full_adder fa_4_39_3(.S(p_4_39[7]), .Cout(p_4_40[3]), .A(p_3_39[3]), .B(p_3_39[2]), .Cin(p_3_39[1]));
full_adder fa_4_40_0(.S(p_4_40[4]), .Cout(p_4_41[0]), .A(p_3_40[12]), .B(p_3_40[11]), .Cin(p_3_40[10]));
full_adder fa_4_40_1(.S(p_4_40[5]), .Cout(p_4_41[1]), .A(p_3_40[9]), .B(p_3_40[8]), .Cin(p_3_40[7]));
full_adder fa_4_40_2(.S(p_4_40[6]), .Cout(p_4_41[2]), .A(p_3_40[6]), .B(p_3_40[5]), .Cin(p_3_40[4]));
full_adder fa_4_40_3(.S(p_4_40[7]), .Cout(p_4_41[3]), .A(p_3_40[3]), .B(p_3_40[2]), .Cin(p_3_40[1]));
full_adder fa_4_41_0(.S(p_4_41[4]), .Cout(p_4_42[0]), .A(p_3_41[12]), .B(p_3_41[11]), .Cin(p_3_41[10]));
full_adder fa_4_41_1(.S(p_4_41[5]), .Cout(p_4_42[1]), .A(p_3_41[9]), .B(p_3_41[8]), .Cin(p_3_41[7]));
full_adder fa_4_41_2(.S(p_4_41[6]), .Cout(p_4_42[2]), .A(p_3_41[6]), .B(p_3_41[5]), .Cin(p_3_41[4]));
full_adder fa_4_41_3(.S(p_4_41[7]), .Cout(p_4_42[3]), .A(p_3_41[3]), .B(p_3_41[2]), .Cin(p_3_41[1]));
full_adder fa_4_42_0(.S(p_4_42[4]), .Cout(p_4_43[0]), .A(p_3_42[12]), .B(p_3_42[11]), .Cin(p_3_42[10]));
full_adder fa_4_42_1(.S(p_4_42[5]), .Cout(p_4_43[1]), .A(p_3_42[9]), .B(p_3_42[8]), .Cin(p_3_42[7]));
full_adder fa_4_42_2(.S(p_4_42[6]), .Cout(p_4_43[2]), .A(p_3_42[6]), .B(p_3_42[5]), .Cin(p_3_42[4]));
full_adder fa_4_42_3(.S(p_4_42[7]), .Cout(p_4_43[3]), .A(p_3_42[3]), .B(p_3_42[2]), .Cin(p_3_42[1]));
full_adder fa_4_43_0(.S(p_4_43[4]), .Cout(p_4_44[0]), .A(p_3_43[12]), .B(p_3_43[11]), .Cin(p_3_43[10]));
full_adder fa_4_43_1(.S(p_4_43[5]), .Cout(p_4_44[1]), .A(p_3_43[9]), .B(p_3_43[8]), .Cin(p_3_43[7]));
full_adder fa_4_43_2(.S(p_4_43[6]), .Cout(p_4_44[2]), .A(p_3_43[6]), .B(p_3_43[5]), .Cin(p_3_43[4]));
full_adder fa_4_43_3(.S(p_4_43[7]), .Cout(p_4_44[3]), .A(p_3_43[3]), .B(p_3_43[2]), .Cin(p_3_43[1]));
full_adder fa_4_44_0(.S(p_4_44[4]), .Cout(p_4_45[0]), .A(p_3_44[12]), .B(p_3_44[11]), .Cin(p_3_44[10]));
full_adder fa_4_44_1(.S(p_4_44[5]), .Cout(p_4_45[1]), .A(p_3_44[9]), .B(p_3_44[8]), .Cin(p_3_44[7]));
full_adder fa_4_44_2(.S(p_4_44[6]), .Cout(p_4_45[2]), .A(p_3_44[6]), .B(p_3_44[5]), .Cin(p_3_44[4]));
full_adder fa_4_44_3(.S(p_4_44[7]), .Cout(p_4_45[3]), .A(p_3_44[3]), .B(p_3_44[2]), .Cin(p_3_44[1]));
full_adder fa_4_45_0(.S(p_4_45[4]), .Cout(p_4_46[0]), .A(p_3_45[12]), .B(p_3_45[11]), .Cin(p_3_45[10]));
full_adder fa_4_45_1(.S(p_4_45[5]), .Cout(p_4_46[1]), .A(p_3_45[9]), .B(p_3_45[8]), .Cin(p_3_45[7]));
full_adder fa_4_45_2(.S(p_4_45[6]), .Cout(p_4_46[2]), .A(p_3_45[6]), .B(p_3_45[5]), .Cin(p_3_45[4]));
full_adder fa_4_45_3(.S(p_4_45[7]), .Cout(p_4_46[3]), .A(p_3_45[3]), .B(p_3_45[2]), .Cin(p_3_45[1]));
full_adder fa_4_46_0(.S(p_4_46[4]), .Cout(p_4_47[0]), .A(p_3_46[12]), .B(p_3_46[11]), .Cin(p_3_46[10]));
full_adder fa_4_46_1(.S(p_4_46[5]), .Cout(p_4_47[1]), .A(p_3_46[9]), .B(p_3_46[8]), .Cin(p_3_46[7]));
full_adder fa_4_46_2(.S(p_4_46[6]), .Cout(p_4_47[2]), .A(p_3_46[6]), .B(p_3_46[5]), .Cin(p_3_46[4]));
full_adder fa_4_46_3(.S(p_4_46[7]), .Cout(p_4_47[3]), .A(p_3_46[3]), .B(p_3_46[2]), .Cin(p_3_46[1]));
full_adder fa_4_47_0(.S(p_4_47[4]), .Cout(p_4_48[0]), .A(p_3_47[12]), .B(p_3_47[11]), .Cin(p_3_47[10]));
full_adder fa_4_47_1(.S(p_4_47[5]), .Cout(p_4_48[1]), .A(p_3_47[9]), .B(p_3_47[8]), .Cin(p_3_47[7]));
full_adder fa_4_47_2(.S(p_4_47[6]), .Cout(p_4_48[2]), .A(p_3_47[6]), .B(p_3_47[5]), .Cin(p_3_47[4]));
full_adder fa_4_47_3(.S(p_4_47[7]), .Cout(p_4_48[3]), .A(p_3_47[3]), .B(p_3_47[2]), .Cin(p_3_47[1]));
full_adder fa_4_48_0(.S(p_4_48[4]), .Cout(p_4_49[0]), .A(p_3_48[12]), .B(p_3_48[11]), .Cin(p_3_48[10]));
full_adder fa_4_48_1(.S(p_4_48[5]), .Cout(p_4_49[1]), .A(p_3_48[9]), .B(p_3_48[8]), .Cin(p_3_48[7]));
full_adder fa_4_48_2(.S(p_4_48[6]), .Cout(p_4_49[2]), .A(p_3_48[6]), .B(p_3_48[5]), .Cin(p_3_48[4]));
full_adder fa_4_48_3(.S(p_4_48[7]), .Cout(p_4_49[3]), .A(p_3_48[3]), .B(p_3_48[2]), .Cin(p_3_48[1]));
full_adder fa_4_49_0(.S(p_4_49[4]), .Cout(p_4_50[0]), .A(p_3_49[12]), .B(p_3_49[11]), .Cin(p_3_49[10]));
full_adder fa_4_49_1(.S(p_4_49[5]), .Cout(p_4_50[1]), .A(p_3_49[9]), .B(p_3_49[8]), .Cin(p_3_49[7]));
full_adder fa_4_49_2(.S(p_4_49[6]), .Cout(p_4_50[2]), .A(p_3_49[6]), .B(p_3_49[5]), .Cin(p_3_49[4]));
full_adder fa_4_49_3(.S(p_4_49[7]), .Cout(p_4_50[3]), .A(p_3_49[3]), .B(p_3_49[2]), .Cin(p_3_49[1]));
full_adder fa_4_50_0(.S(p_4_50[4]), .Cout(p_4_51[0]), .A(p_3_50[12]), .B(p_3_50[11]), .Cin(p_3_50[10]));
full_adder fa_4_50_1(.S(p_4_50[5]), .Cout(p_4_51[1]), .A(p_3_50[9]), .B(p_3_50[8]), .Cin(p_3_50[7]));
full_adder fa_4_50_2(.S(p_4_50[6]), .Cout(p_4_51[2]), .A(p_3_50[6]), .B(p_3_50[5]), .Cin(p_3_50[4]));
full_adder fa_4_50_3(.S(p_4_50[7]), .Cout(p_4_51[3]), .A(p_3_50[3]), .B(p_3_50[2]), .Cin(p_3_50[1]));
full_adder fa_4_51_0(.S(p_4_51[4]), .Cout(p_4_52[0]), .A(p_3_51[12]), .B(p_3_51[11]), .Cin(p_3_51[10]));
full_adder fa_4_51_1(.S(p_4_51[5]), .Cout(p_4_52[1]), .A(p_3_51[9]), .B(p_3_51[8]), .Cin(p_3_51[7]));
full_adder fa_4_51_2(.S(p_4_51[6]), .Cout(p_4_52[2]), .A(p_3_51[6]), .B(p_3_51[5]), .Cin(p_3_51[4]));
full_adder fa_4_51_3(.S(p_4_51[7]), .Cout(p_4_52[3]), .A(p_3_51[3]), .B(p_3_51[2]), .Cin(p_3_51[1]));
full_adder fa_4_52_0(.S(p_4_52[4]), .Cout(p_4_53[0]), .A(p_3_52[10]), .B(p_3_52[9]), .Cin(p_3_52[8]));
full_adder fa_4_52_1(.S(p_4_52[5]), .Cout(p_4_53[1]), .A(p_3_52[7]), .B(p_3_52[6]), .Cin(p_3_52[5]));
full_adder fa_4_52_2(.S(p_4_52[6]), .Cout(p_4_53[2]), .A(p_3_52[4]), .B(p_3_52[3]), .Cin(p_3_52[2]));
full_adder fa_4_53_0(.S(p_4_53[3]), .Cout(p_4_54[0]), .A(p_3_53[9]), .B(p_3_53[8]), .Cin(p_3_53[7]));
full_adder fa_4_53_1(.S(p_4_53[4]), .Cout(p_4_54[1]), .A(p_3_53[6]), .B(p_3_53[5]), .Cin(p_3_53[4]));
full_adder fa_4_54_0(.S(p_4_54[2]), .Cout(p_4_55[0]), .A(p_3_54[8]), .B(p_3_54[7]), .Cin(p_3_54[6]));

// Stage 5 non-added partial products
assign p_5_0[0:0] = p_4_0[0:0];
assign p_5_1[1:0] = p_4_1[1:0];
assign p_5_2[2:0] = p_4_2[2:0];
assign p_5_3[3:0] = p_4_3[3:0];
assign p_5_4[4:0] = p_4_4[4:0];
assign p_5_5[5:0] = p_4_5[5:0];
assign p_5_6[5:1] = p_4_6[4:0];
assign p_5_7[5:3] = p_4_7[2:0];
assign p_5_8[5:5] = p_4_8[0:0];
assign p_5_56[5:5] = p_4_56[0:0];
assign p_5_57[5:3] = p_4_57[2:0];
assign p_5_58[5:1] = p_4_58[4:0];
assign p_5_59[3:0] = p_4_59[3:0];
assign p_5_60[2:0] = p_4_60[2:0];
assign p_5_61[1:0] = p_4_61[1:0];
assign p_5_62[0:0] = p_4_62[0:0];
// Stage 5 adders
half_adder ha_5_6(.S(p_5_6[0]), .Cout(p_5_7[0]), .A(p_4_6[6]), .B(p_4_6[5]));
full_adder fa_5_7_0(.S(p_5_7[1]), .Cout(p_5_8[0]), .A(p_4_7[7]), .B(p_4_7[6]), .Cin(p_4_7[5]));
half_adder ha_5_7(.S(p_5_7[2]), .Cout(p_5_8[1]), .A(p_4_7[4]), .B(p_4_7[3]));
full_adder fa_5_8_0(.S(p_5_8[2]), .Cout(p_5_9[0]), .A(p_4_8[8]), .B(p_4_8[7]), .Cin(p_4_8[6]));
full_adder fa_5_8_1(.S(p_5_8[3]), .Cout(p_5_9[1]), .A(p_4_8[5]), .B(p_4_8[4]), .Cin(p_4_8[3]));
half_adder ha_5_8(.S(p_5_8[4]), .Cout(p_5_9[2]), .A(p_4_8[2]), .B(p_4_8[1]));
full_adder fa_5_9_0(.S(p_5_9[3]), .Cout(p_5_10[0]), .A(p_4_9[8]), .B(p_4_9[7]), .Cin(p_4_9[6]));
full_adder fa_5_9_1(.S(p_5_9[4]), .Cout(p_5_10[1]), .A(p_4_9[5]), .B(p_4_9[4]), .Cin(p_4_9[3]));
full_adder fa_5_9_2(.S(p_5_9[5]), .Cout(p_5_10[2]), .A(p_4_9[2]), .B(p_4_9[1]), .Cin(p_4_9[0]));
full_adder fa_5_10_0(.S(p_5_10[3]), .Cout(p_5_11[0]), .A(p_4_10[8]), .B(p_4_10[7]), .Cin(p_4_10[6]));
full_adder fa_5_10_1(.S(p_5_10[4]), .Cout(p_5_11[1]), .A(p_4_10[5]), .B(p_4_10[4]), .Cin(p_4_10[3]));
full_adder fa_5_10_2(.S(p_5_10[5]), .Cout(p_5_11[2]), .A(p_4_10[2]), .B(p_4_10[1]), .Cin(p_4_10[0]));
full_adder fa_5_11_0(.S(p_5_11[3]), .Cout(p_5_12[0]), .A(p_4_11[8]), .B(p_4_11[7]), .Cin(p_4_11[6]));
full_adder fa_5_11_1(.S(p_5_11[4]), .Cout(p_5_12[1]), .A(p_4_11[5]), .B(p_4_11[4]), .Cin(p_4_11[3]));
full_adder fa_5_11_2(.S(p_5_11[5]), .Cout(p_5_12[2]), .A(p_4_11[2]), .B(p_4_11[1]), .Cin(p_4_11[0]));
full_adder fa_5_12_0(.S(p_5_12[3]), .Cout(p_5_13[0]), .A(p_4_12[8]), .B(p_4_12[7]), .Cin(p_4_12[6]));
full_adder fa_5_12_1(.S(p_5_12[4]), .Cout(p_5_13[1]), .A(p_4_12[5]), .B(p_4_12[4]), .Cin(p_4_12[3]));
full_adder fa_5_12_2(.S(p_5_12[5]), .Cout(p_5_13[2]), .A(p_4_12[2]), .B(p_4_12[1]), .Cin(p_4_12[0]));
full_adder fa_5_13_0(.S(p_5_13[3]), .Cout(p_5_14[0]), .A(p_4_13[8]), .B(p_4_13[7]), .Cin(p_4_13[6]));
full_adder fa_5_13_1(.S(p_5_13[4]), .Cout(p_5_14[1]), .A(p_4_13[5]), .B(p_4_13[4]), .Cin(p_4_13[3]));
full_adder fa_5_13_2(.S(p_5_13[5]), .Cout(p_5_14[2]), .A(p_4_13[2]), .B(p_4_13[1]), .Cin(p_4_13[0]));
full_adder fa_5_14_0(.S(p_5_14[3]), .Cout(p_5_15[0]), .A(p_4_14[8]), .B(p_4_14[7]), .Cin(p_4_14[6]));
full_adder fa_5_14_1(.S(p_5_14[4]), .Cout(p_5_15[1]), .A(p_4_14[5]), .B(p_4_14[4]), .Cin(p_4_14[3]));
full_adder fa_5_14_2(.S(p_5_14[5]), .Cout(p_5_15[2]), .A(p_4_14[2]), .B(p_4_14[1]), .Cin(p_4_14[0]));
full_adder fa_5_15_0(.S(p_5_15[3]), .Cout(p_5_16[0]), .A(p_4_15[8]), .B(p_4_15[7]), .Cin(p_4_15[6]));
full_adder fa_5_15_1(.S(p_5_15[4]), .Cout(p_5_16[1]), .A(p_4_15[5]), .B(p_4_15[4]), .Cin(p_4_15[3]));
full_adder fa_5_15_2(.S(p_5_15[5]), .Cout(p_5_16[2]), .A(p_4_15[2]), .B(p_4_15[1]), .Cin(p_4_15[0]));
full_adder fa_5_16_0(.S(p_5_16[3]), .Cout(p_5_17[0]), .A(p_4_16[8]), .B(p_4_16[7]), .Cin(p_4_16[6]));
full_adder fa_5_16_1(.S(p_5_16[4]), .Cout(p_5_17[1]), .A(p_4_16[5]), .B(p_4_16[4]), .Cin(p_4_16[3]));
full_adder fa_5_16_2(.S(p_5_16[5]), .Cout(p_5_17[2]), .A(p_4_16[2]), .B(p_4_16[1]), .Cin(p_4_16[0]));
full_adder fa_5_17_0(.S(p_5_17[3]), .Cout(p_5_18[0]), .A(p_4_17[8]), .B(p_4_17[7]), .Cin(p_4_17[6]));
full_adder fa_5_17_1(.S(p_5_17[4]), .Cout(p_5_18[1]), .A(p_4_17[5]), .B(p_4_17[4]), .Cin(p_4_17[3]));
full_adder fa_5_17_2(.S(p_5_17[5]), .Cout(p_5_18[2]), .A(p_4_17[2]), .B(p_4_17[1]), .Cin(p_4_17[0]));
full_adder fa_5_18_0(.S(p_5_18[3]), .Cout(p_5_19[0]), .A(p_4_18[8]), .B(p_4_18[7]), .Cin(p_4_18[6]));
full_adder fa_5_18_1(.S(p_5_18[4]), .Cout(p_5_19[1]), .A(p_4_18[5]), .B(p_4_18[4]), .Cin(p_4_18[3]));
full_adder fa_5_18_2(.S(p_5_18[5]), .Cout(p_5_19[2]), .A(p_4_18[2]), .B(p_4_18[1]), .Cin(p_4_18[0]));
full_adder fa_5_19_0(.S(p_5_19[3]), .Cout(p_5_20[0]), .A(p_4_19[8]), .B(p_4_19[7]), .Cin(p_4_19[6]));
full_adder fa_5_19_1(.S(p_5_19[4]), .Cout(p_5_20[1]), .A(p_4_19[5]), .B(p_4_19[4]), .Cin(p_4_19[3]));
full_adder fa_5_19_2(.S(p_5_19[5]), .Cout(p_5_20[2]), .A(p_4_19[2]), .B(p_4_19[1]), .Cin(p_4_19[0]));
full_adder fa_5_20_0(.S(p_5_20[3]), .Cout(p_5_21[0]), .A(p_4_20[8]), .B(p_4_20[7]), .Cin(p_4_20[6]));
full_adder fa_5_20_1(.S(p_5_20[4]), .Cout(p_5_21[1]), .A(p_4_20[5]), .B(p_4_20[4]), .Cin(p_4_20[3]));
full_adder fa_5_20_2(.S(p_5_20[5]), .Cout(p_5_21[2]), .A(p_4_20[2]), .B(p_4_20[1]), .Cin(p_4_20[0]));
full_adder fa_5_21_0(.S(p_5_21[3]), .Cout(p_5_22[0]), .A(p_4_21[8]), .B(p_4_21[7]), .Cin(p_4_21[6]));
full_adder fa_5_21_1(.S(p_5_21[4]), .Cout(p_5_22[1]), .A(p_4_21[5]), .B(p_4_21[4]), .Cin(p_4_21[3]));
full_adder fa_5_21_2(.S(p_5_21[5]), .Cout(p_5_22[2]), .A(p_4_21[2]), .B(p_4_21[1]), .Cin(p_4_21[0]));
full_adder fa_5_22_0(.S(p_5_22[3]), .Cout(p_5_23[0]), .A(p_4_22[8]), .B(p_4_22[7]), .Cin(p_4_22[6]));
full_adder fa_5_22_1(.S(p_5_22[4]), .Cout(p_5_23[1]), .A(p_4_22[5]), .B(p_4_22[4]), .Cin(p_4_22[3]));
full_adder fa_5_22_2(.S(p_5_22[5]), .Cout(p_5_23[2]), .A(p_4_22[2]), .B(p_4_22[1]), .Cin(p_4_22[0]));
full_adder fa_5_23_0(.S(p_5_23[3]), .Cout(p_5_24[0]), .A(p_4_23[8]), .B(p_4_23[7]), .Cin(p_4_23[6]));
full_adder fa_5_23_1(.S(p_5_23[4]), .Cout(p_5_24[1]), .A(p_4_23[5]), .B(p_4_23[4]), .Cin(p_4_23[3]));
full_adder fa_5_23_2(.S(p_5_23[5]), .Cout(p_5_24[2]), .A(p_4_23[2]), .B(p_4_23[1]), .Cin(p_4_23[0]));
full_adder fa_5_24_0(.S(p_5_24[3]), .Cout(p_5_25[0]), .A(p_4_24[8]), .B(p_4_24[7]), .Cin(p_4_24[6]));
full_adder fa_5_24_1(.S(p_5_24[4]), .Cout(p_5_25[1]), .A(p_4_24[5]), .B(p_4_24[4]), .Cin(p_4_24[3]));
full_adder fa_5_24_2(.S(p_5_24[5]), .Cout(p_5_25[2]), .A(p_4_24[2]), .B(p_4_24[1]), .Cin(p_4_24[0]));
full_adder fa_5_25_0(.S(p_5_25[3]), .Cout(p_5_26[0]), .A(p_4_25[8]), .B(p_4_25[7]), .Cin(p_4_25[6]));
full_adder fa_5_25_1(.S(p_5_25[4]), .Cout(p_5_26[1]), .A(p_4_25[5]), .B(p_4_25[4]), .Cin(p_4_25[3]));
full_adder fa_5_25_2(.S(p_5_25[5]), .Cout(p_5_26[2]), .A(p_4_25[2]), .B(p_4_25[1]), .Cin(p_4_25[0]));
full_adder fa_5_26_0(.S(p_5_26[3]), .Cout(p_5_27[0]), .A(p_4_26[8]), .B(p_4_26[7]), .Cin(p_4_26[6]));
full_adder fa_5_26_1(.S(p_5_26[4]), .Cout(p_5_27[1]), .A(p_4_26[5]), .B(p_4_26[4]), .Cin(p_4_26[3]));
full_adder fa_5_26_2(.S(p_5_26[5]), .Cout(p_5_27[2]), .A(p_4_26[2]), .B(p_4_26[1]), .Cin(p_4_26[0]));
full_adder fa_5_27_0(.S(p_5_27[3]), .Cout(p_5_28[0]), .A(p_4_27[8]), .B(p_4_27[7]), .Cin(p_4_27[6]));
full_adder fa_5_27_1(.S(p_5_27[4]), .Cout(p_5_28[1]), .A(p_4_27[5]), .B(p_4_27[4]), .Cin(p_4_27[3]));
full_adder fa_5_27_2(.S(p_5_27[5]), .Cout(p_5_28[2]), .A(p_4_27[2]), .B(p_4_27[1]), .Cin(p_4_27[0]));
full_adder fa_5_28_0(.S(p_5_28[3]), .Cout(p_5_29[0]), .A(p_4_28[8]), .B(p_4_28[7]), .Cin(p_4_28[6]));
full_adder fa_5_28_1(.S(p_5_28[4]), .Cout(p_5_29[1]), .A(p_4_28[5]), .B(p_4_28[4]), .Cin(p_4_28[3]));
full_adder fa_5_28_2(.S(p_5_28[5]), .Cout(p_5_29[2]), .A(p_4_28[2]), .B(p_4_28[1]), .Cin(p_4_28[0]));
full_adder fa_5_29_0(.S(p_5_29[3]), .Cout(p_5_30[0]), .A(p_4_29[8]), .B(p_4_29[7]), .Cin(p_4_29[6]));
full_adder fa_5_29_1(.S(p_5_29[4]), .Cout(p_5_30[1]), .A(p_4_29[5]), .B(p_4_29[4]), .Cin(p_4_29[3]));
full_adder fa_5_29_2(.S(p_5_29[5]), .Cout(p_5_30[2]), .A(p_4_29[2]), .B(p_4_29[1]), .Cin(p_4_29[0]));
full_adder fa_5_30_0(.S(p_5_30[3]), .Cout(p_5_31[0]), .A(p_4_30[8]), .B(p_4_30[7]), .Cin(p_4_30[6]));
full_adder fa_5_30_1(.S(p_5_30[4]), .Cout(p_5_31[1]), .A(p_4_30[5]), .B(p_4_30[4]), .Cin(p_4_30[3]));
full_adder fa_5_30_2(.S(p_5_30[5]), .Cout(p_5_31[2]), .A(p_4_30[2]), .B(p_4_30[1]), .Cin(p_4_30[0]));
full_adder fa_5_31_0(.S(p_5_31[3]), .Cout(p_5_32[0]), .A(p_4_31[8]), .B(p_4_31[7]), .Cin(p_4_31[6]));
full_adder fa_5_31_1(.S(p_5_31[4]), .Cout(p_5_32[1]), .A(p_4_31[5]), .B(p_4_31[4]), .Cin(p_4_31[3]));
full_adder fa_5_31_2(.S(p_5_31[5]), .Cout(p_5_32[2]), .A(p_4_31[2]), .B(p_4_31[1]), .Cin(p_4_31[0]));
full_adder fa_5_32_0(.S(p_5_32[3]), .Cout(p_5_33[0]), .A(p_4_32[8]), .B(p_4_32[7]), .Cin(p_4_32[6]));
full_adder fa_5_32_1(.S(p_5_32[4]), .Cout(p_5_33[1]), .A(p_4_32[5]), .B(p_4_32[4]), .Cin(p_4_32[3]));
full_adder fa_5_32_2(.S(p_5_32[5]), .Cout(p_5_33[2]), .A(p_4_32[2]), .B(p_4_32[1]), .Cin(p_4_32[0]));
full_adder fa_5_33_0(.S(p_5_33[3]), .Cout(p_5_34[0]), .A(p_4_33[8]), .B(p_4_33[7]), .Cin(p_4_33[6]));
full_adder fa_5_33_1(.S(p_5_33[4]), .Cout(p_5_34[1]), .A(p_4_33[5]), .B(p_4_33[4]), .Cin(p_4_33[3]));
full_adder fa_5_33_2(.S(p_5_33[5]), .Cout(p_5_34[2]), .A(p_4_33[2]), .B(p_4_33[1]), .Cin(p_4_33[0]));
full_adder fa_5_34_0(.S(p_5_34[3]), .Cout(p_5_35[0]), .A(p_4_34[8]), .B(p_4_34[7]), .Cin(p_4_34[6]));
full_adder fa_5_34_1(.S(p_5_34[4]), .Cout(p_5_35[1]), .A(p_4_34[5]), .B(p_4_34[4]), .Cin(p_4_34[3]));
full_adder fa_5_34_2(.S(p_5_34[5]), .Cout(p_5_35[2]), .A(p_4_34[2]), .B(p_4_34[1]), .Cin(p_4_34[0]));
full_adder fa_5_35_0(.S(p_5_35[3]), .Cout(p_5_36[0]), .A(p_4_35[8]), .B(p_4_35[7]), .Cin(p_4_35[6]));
full_adder fa_5_35_1(.S(p_5_35[4]), .Cout(p_5_36[1]), .A(p_4_35[5]), .B(p_4_35[4]), .Cin(p_4_35[3]));
full_adder fa_5_35_2(.S(p_5_35[5]), .Cout(p_5_36[2]), .A(p_4_35[2]), .B(p_4_35[1]), .Cin(p_4_35[0]));
full_adder fa_5_36_0(.S(p_5_36[3]), .Cout(p_5_37[0]), .A(p_4_36[8]), .B(p_4_36[7]), .Cin(p_4_36[6]));
full_adder fa_5_36_1(.S(p_5_36[4]), .Cout(p_5_37[1]), .A(p_4_36[5]), .B(p_4_36[4]), .Cin(p_4_36[3]));
full_adder fa_5_36_2(.S(p_5_36[5]), .Cout(p_5_37[2]), .A(p_4_36[2]), .B(p_4_36[1]), .Cin(p_4_36[0]));
full_adder fa_5_37_0(.S(p_5_37[3]), .Cout(p_5_38[0]), .A(p_4_37[8]), .B(p_4_37[7]), .Cin(p_4_37[6]));
full_adder fa_5_37_1(.S(p_5_37[4]), .Cout(p_5_38[1]), .A(p_4_37[5]), .B(p_4_37[4]), .Cin(p_4_37[3]));
full_adder fa_5_37_2(.S(p_5_37[5]), .Cout(p_5_38[2]), .A(p_4_37[2]), .B(p_4_37[1]), .Cin(p_4_37[0]));
full_adder fa_5_38_0(.S(p_5_38[3]), .Cout(p_5_39[0]), .A(p_4_38[8]), .B(p_4_38[7]), .Cin(p_4_38[6]));
full_adder fa_5_38_1(.S(p_5_38[4]), .Cout(p_5_39[1]), .A(p_4_38[5]), .B(p_4_38[4]), .Cin(p_4_38[3]));
full_adder fa_5_38_2(.S(p_5_38[5]), .Cout(p_5_39[2]), .A(p_4_38[2]), .B(p_4_38[1]), .Cin(p_4_38[0]));
full_adder fa_5_39_0(.S(p_5_39[3]), .Cout(p_5_40[0]), .A(p_4_39[8]), .B(p_4_39[7]), .Cin(p_4_39[6]));
full_adder fa_5_39_1(.S(p_5_39[4]), .Cout(p_5_40[1]), .A(p_4_39[5]), .B(p_4_39[4]), .Cin(p_4_39[3]));
full_adder fa_5_39_2(.S(p_5_39[5]), .Cout(p_5_40[2]), .A(p_4_39[2]), .B(p_4_39[1]), .Cin(p_4_39[0]));
full_adder fa_5_40_0(.S(p_5_40[3]), .Cout(p_5_41[0]), .A(p_4_40[8]), .B(p_4_40[7]), .Cin(p_4_40[6]));
full_adder fa_5_40_1(.S(p_5_40[4]), .Cout(p_5_41[1]), .A(p_4_40[5]), .B(p_4_40[4]), .Cin(p_4_40[3]));
full_adder fa_5_40_2(.S(p_5_40[5]), .Cout(p_5_41[2]), .A(p_4_40[2]), .B(p_4_40[1]), .Cin(p_4_40[0]));
full_adder fa_5_41_0(.S(p_5_41[3]), .Cout(p_5_42[0]), .A(p_4_41[8]), .B(p_4_41[7]), .Cin(p_4_41[6]));
full_adder fa_5_41_1(.S(p_5_41[4]), .Cout(p_5_42[1]), .A(p_4_41[5]), .B(p_4_41[4]), .Cin(p_4_41[3]));
full_adder fa_5_41_2(.S(p_5_41[5]), .Cout(p_5_42[2]), .A(p_4_41[2]), .B(p_4_41[1]), .Cin(p_4_41[0]));
full_adder fa_5_42_0(.S(p_5_42[3]), .Cout(p_5_43[0]), .A(p_4_42[8]), .B(p_4_42[7]), .Cin(p_4_42[6]));
full_adder fa_5_42_1(.S(p_5_42[4]), .Cout(p_5_43[1]), .A(p_4_42[5]), .B(p_4_42[4]), .Cin(p_4_42[3]));
full_adder fa_5_42_2(.S(p_5_42[5]), .Cout(p_5_43[2]), .A(p_4_42[2]), .B(p_4_42[1]), .Cin(p_4_42[0]));
full_adder fa_5_43_0(.S(p_5_43[3]), .Cout(p_5_44[0]), .A(p_4_43[8]), .B(p_4_43[7]), .Cin(p_4_43[6]));
full_adder fa_5_43_1(.S(p_5_43[4]), .Cout(p_5_44[1]), .A(p_4_43[5]), .B(p_4_43[4]), .Cin(p_4_43[3]));
full_adder fa_5_43_2(.S(p_5_43[5]), .Cout(p_5_44[2]), .A(p_4_43[2]), .B(p_4_43[1]), .Cin(p_4_43[0]));
full_adder fa_5_44_0(.S(p_5_44[3]), .Cout(p_5_45[0]), .A(p_4_44[8]), .B(p_4_44[7]), .Cin(p_4_44[6]));
full_adder fa_5_44_1(.S(p_5_44[4]), .Cout(p_5_45[1]), .A(p_4_44[5]), .B(p_4_44[4]), .Cin(p_4_44[3]));
full_adder fa_5_44_2(.S(p_5_44[5]), .Cout(p_5_45[2]), .A(p_4_44[2]), .B(p_4_44[1]), .Cin(p_4_44[0]));
full_adder fa_5_45_0(.S(p_5_45[3]), .Cout(p_5_46[0]), .A(p_4_45[8]), .B(p_4_45[7]), .Cin(p_4_45[6]));
full_adder fa_5_45_1(.S(p_5_45[4]), .Cout(p_5_46[1]), .A(p_4_45[5]), .B(p_4_45[4]), .Cin(p_4_45[3]));
full_adder fa_5_45_2(.S(p_5_45[5]), .Cout(p_5_46[2]), .A(p_4_45[2]), .B(p_4_45[1]), .Cin(p_4_45[0]));
full_adder fa_5_46_0(.S(p_5_46[3]), .Cout(p_5_47[0]), .A(p_4_46[8]), .B(p_4_46[7]), .Cin(p_4_46[6]));
full_adder fa_5_46_1(.S(p_5_46[4]), .Cout(p_5_47[1]), .A(p_4_46[5]), .B(p_4_46[4]), .Cin(p_4_46[3]));
full_adder fa_5_46_2(.S(p_5_46[5]), .Cout(p_5_47[2]), .A(p_4_46[2]), .B(p_4_46[1]), .Cin(p_4_46[0]));
full_adder fa_5_47_0(.S(p_5_47[3]), .Cout(p_5_48[0]), .A(p_4_47[8]), .B(p_4_47[7]), .Cin(p_4_47[6]));
full_adder fa_5_47_1(.S(p_5_47[4]), .Cout(p_5_48[1]), .A(p_4_47[5]), .B(p_4_47[4]), .Cin(p_4_47[3]));
full_adder fa_5_47_2(.S(p_5_47[5]), .Cout(p_5_48[2]), .A(p_4_47[2]), .B(p_4_47[1]), .Cin(p_4_47[0]));
full_adder fa_5_48_0(.S(p_5_48[3]), .Cout(p_5_49[0]), .A(p_4_48[8]), .B(p_4_48[7]), .Cin(p_4_48[6]));
full_adder fa_5_48_1(.S(p_5_48[4]), .Cout(p_5_49[1]), .A(p_4_48[5]), .B(p_4_48[4]), .Cin(p_4_48[3]));
full_adder fa_5_48_2(.S(p_5_48[5]), .Cout(p_5_49[2]), .A(p_4_48[2]), .B(p_4_48[1]), .Cin(p_4_48[0]));
full_adder fa_5_49_0(.S(p_5_49[3]), .Cout(p_5_50[0]), .A(p_4_49[8]), .B(p_4_49[7]), .Cin(p_4_49[6]));
full_adder fa_5_49_1(.S(p_5_49[4]), .Cout(p_5_50[1]), .A(p_4_49[5]), .B(p_4_49[4]), .Cin(p_4_49[3]));
full_adder fa_5_49_2(.S(p_5_49[5]), .Cout(p_5_50[2]), .A(p_4_49[2]), .B(p_4_49[1]), .Cin(p_4_49[0]));
full_adder fa_5_50_0(.S(p_5_50[3]), .Cout(p_5_51[0]), .A(p_4_50[8]), .B(p_4_50[7]), .Cin(p_4_50[6]));
full_adder fa_5_50_1(.S(p_5_50[4]), .Cout(p_5_51[1]), .A(p_4_50[5]), .B(p_4_50[4]), .Cin(p_4_50[3]));
full_adder fa_5_50_2(.S(p_5_50[5]), .Cout(p_5_51[2]), .A(p_4_50[2]), .B(p_4_50[1]), .Cin(p_4_50[0]));
full_adder fa_5_51_0(.S(p_5_51[3]), .Cout(p_5_52[0]), .A(p_4_51[8]), .B(p_4_51[7]), .Cin(p_4_51[6]));
full_adder fa_5_51_1(.S(p_5_51[4]), .Cout(p_5_52[1]), .A(p_4_51[5]), .B(p_4_51[4]), .Cin(p_4_51[3]));
full_adder fa_5_51_2(.S(p_5_51[5]), .Cout(p_5_52[2]), .A(p_4_51[2]), .B(p_4_51[1]), .Cin(p_4_51[0]));
full_adder fa_5_52_0(.S(p_5_52[3]), .Cout(p_5_53[0]), .A(p_4_52[8]), .B(p_4_52[7]), .Cin(p_4_52[6]));
full_adder fa_5_52_1(.S(p_5_52[4]), .Cout(p_5_53[1]), .A(p_4_52[5]), .B(p_4_52[4]), .Cin(p_4_52[3]));
full_adder fa_5_52_2(.S(p_5_52[5]), .Cout(p_5_53[2]), .A(p_4_52[2]), .B(p_4_52[1]), .Cin(p_4_52[0]));
full_adder fa_5_53_0(.S(p_5_53[3]), .Cout(p_5_54[0]), .A(p_4_53[8]), .B(p_4_53[7]), .Cin(p_4_53[6]));
full_adder fa_5_53_1(.S(p_5_53[4]), .Cout(p_5_54[1]), .A(p_4_53[5]), .B(p_4_53[4]), .Cin(p_4_53[3]));
full_adder fa_5_53_2(.S(p_5_53[5]), .Cout(p_5_54[2]), .A(p_4_53[2]), .B(p_4_53[1]), .Cin(p_4_53[0]));
full_adder fa_5_54_0(.S(p_5_54[3]), .Cout(p_5_55[0]), .A(p_4_54[8]), .B(p_4_54[7]), .Cin(p_4_54[6]));
full_adder fa_5_54_1(.S(p_5_54[4]), .Cout(p_5_55[1]), .A(p_4_54[5]), .B(p_4_54[4]), .Cin(p_4_54[3]));
full_adder fa_5_54_2(.S(p_5_54[5]), .Cout(p_5_55[2]), .A(p_4_54[2]), .B(p_4_54[1]), .Cin(p_4_54[0]));
full_adder fa_5_55_0(.S(p_5_55[3]), .Cout(p_5_56[0]), .A(p_4_55[8]), .B(p_4_55[7]), .Cin(p_4_55[6]));
full_adder fa_5_55_1(.S(p_5_55[4]), .Cout(p_5_56[1]), .A(p_4_55[5]), .B(p_4_55[4]), .Cin(p_4_55[3]));
full_adder fa_5_55_2(.S(p_5_55[5]), .Cout(p_5_56[2]), .A(p_4_55[2]), .B(p_4_55[1]), .Cin(p_4_55[0]));
full_adder fa_5_56_0(.S(p_5_56[3]), .Cout(p_5_57[0]), .A(p_4_56[6]), .B(p_4_56[5]), .Cin(p_4_56[4]));
full_adder fa_5_56_1(.S(p_5_56[4]), .Cout(p_5_57[1]), .A(p_4_56[3]), .B(p_4_56[2]), .Cin(p_4_56[1]));
full_adder fa_5_57_0(.S(p_5_57[2]), .Cout(p_5_58[0]), .A(p_4_57[5]), .B(p_4_57[4]), .Cin(p_4_57[3]));

// Stage 6 non-added partial products
assign p_6_0[0:0] = p_5_0[0:0];
assign p_6_1[1:0] = p_5_1[1:0];
assign p_6_2[2:0] = p_5_2[2:0];
assign p_6_3[3:0] = p_5_3[3:0];
assign p_6_4[3:1] = p_5_4[2:0];
assign p_6_5[3:3] = p_5_5[0:0];
assign p_6_59[3:3] = p_5_59[0:0];
assign p_6_60[3:1] = p_5_60[2:0];
assign p_6_61[1:0] = p_5_61[1:0];
assign p_6_62[0:0] = p_5_62[0:0];
// Stage 6 adders
half_adder ha_6_4(.S(p_6_4[0]), .Cout(p_6_5[0]), .A(p_5_4[4]), .B(p_5_4[3]));
full_adder fa_6_5_0(.S(p_6_5[1]), .Cout(p_6_6[0]), .A(p_5_5[5]), .B(p_5_5[4]), .Cin(p_5_5[3]));
half_adder ha_6_5(.S(p_6_5[2]), .Cout(p_6_6[1]), .A(p_5_5[2]), .B(p_5_5[1]));
full_adder fa_6_6_0(.S(p_6_6[2]), .Cout(p_6_7[0]), .A(p_5_6[5]), .B(p_5_6[4]), .Cin(p_5_6[3]));
full_adder fa_6_6_1(.S(p_6_6[3]), .Cout(p_6_7[1]), .A(p_5_6[2]), .B(p_5_6[1]), .Cin(p_5_6[0]));
full_adder fa_6_7_0(.S(p_6_7[2]), .Cout(p_6_8[0]), .A(p_5_7[5]), .B(p_5_7[4]), .Cin(p_5_7[3]));
full_adder fa_6_7_1(.S(p_6_7[3]), .Cout(p_6_8[1]), .A(p_5_7[2]), .B(p_5_7[1]), .Cin(p_5_7[0]));
full_adder fa_6_8_0(.S(p_6_8[2]), .Cout(p_6_9[0]), .A(p_5_8[5]), .B(p_5_8[4]), .Cin(p_5_8[3]));
full_adder fa_6_8_1(.S(p_6_8[3]), .Cout(p_6_9[1]), .A(p_5_8[2]), .B(p_5_8[1]), .Cin(p_5_8[0]));
full_adder fa_6_9_0(.S(p_6_9[2]), .Cout(p_6_10[0]), .A(p_5_9[5]), .B(p_5_9[4]), .Cin(p_5_9[3]));
full_adder fa_6_9_1(.S(p_6_9[3]), .Cout(p_6_10[1]), .A(p_5_9[2]), .B(p_5_9[1]), .Cin(p_5_9[0]));
full_adder fa_6_10_0(.S(p_6_10[2]), .Cout(p_6_11[0]), .A(p_5_10[5]), .B(p_5_10[4]), .Cin(p_5_10[3]));
full_adder fa_6_10_1(.S(p_6_10[3]), .Cout(p_6_11[1]), .A(p_5_10[2]), .B(p_5_10[1]), .Cin(p_5_10[0]));
full_adder fa_6_11_0(.S(p_6_11[2]), .Cout(p_6_12[0]), .A(p_5_11[5]), .B(p_5_11[4]), .Cin(p_5_11[3]));
full_adder fa_6_11_1(.S(p_6_11[3]), .Cout(p_6_12[1]), .A(p_5_11[2]), .B(p_5_11[1]), .Cin(p_5_11[0]));
full_adder fa_6_12_0(.S(p_6_12[2]), .Cout(p_6_13[0]), .A(p_5_12[5]), .B(p_5_12[4]), .Cin(p_5_12[3]));
full_adder fa_6_12_1(.S(p_6_12[3]), .Cout(p_6_13[1]), .A(p_5_12[2]), .B(p_5_12[1]), .Cin(p_5_12[0]));
full_adder fa_6_13_0(.S(p_6_13[2]), .Cout(p_6_14[0]), .A(p_5_13[5]), .B(p_5_13[4]), .Cin(p_5_13[3]));
full_adder fa_6_13_1(.S(p_6_13[3]), .Cout(p_6_14[1]), .A(p_5_13[2]), .B(p_5_13[1]), .Cin(p_5_13[0]));
full_adder fa_6_14_0(.S(p_6_14[2]), .Cout(p_6_15[0]), .A(p_5_14[5]), .B(p_5_14[4]), .Cin(p_5_14[3]));
full_adder fa_6_14_1(.S(p_6_14[3]), .Cout(p_6_15[1]), .A(p_5_14[2]), .B(p_5_14[1]), .Cin(p_5_14[0]));
full_adder fa_6_15_0(.S(p_6_15[2]), .Cout(p_6_16[0]), .A(p_5_15[5]), .B(p_5_15[4]), .Cin(p_5_15[3]));
full_adder fa_6_15_1(.S(p_6_15[3]), .Cout(p_6_16[1]), .A(p_5_15[2]), .B(p_5_15[1]), .Cin(p_5_15[0]));
full_adder fa_6_16_0(.S(p_6_16[2]), .Cout(p_6_17[0]), .A(p_5_16[5]), .B(p_5_16[4]), .Cin(p_5_16[3]));
full_adder fa_6_16_1(.S(p_6_16[3]), .Cout(p_6_17[1]), .A(p_5_16[2]), .B(p_5_16[1]), .Cin(p_5_16[0]));
full_adder fa_6_17_0(.S(p_6_17[2]), .Cout(p_6_18[0]), .A(p_5_17[5]), .B(p_5_17[4]), .Cin(p_5_17[3]));
full_adder fa_6_17_1(.S(p_6_17[3]), .Cout(p_6_18[1]), .A(p_5_17[2]), .B(p_5_17[1]), .Cin(p_5_17[0]));
full_adder fa_6_18_0(.S(p_6_18[2]), .Cout(p_6_19[0]), .A(p_5_18[5]), .B(p_5_18[4]), .Cin(p_5_18[3]));
full_adder fa_6_18_1(.S(p_6_18[3]), .Cout(p_6_19[1]), .A(p_5_18[2]), .B(p_5_18[1]), .Cin(p_5_18[0]));
full_adder fa_6_19_0(.S(p_6_19[2]), .Cout(p_6_20[0]), .A(p_5_19[5]), .B(p_5_19[4]), .Cin(p_5_19[3]));
full_adder fa_6_19_1(.S(p_6_19[3]), .Cout(p_6_20[1]), .A(p_5_19[2]), .B(p_5_19[1]), .Cin(p_5_19[0]));
full_adder fa_6_20_0(.S(p_6_20[2]), .Cout(p_6_21[0]), .A(p_5_20[5]), .B(p_5_20[4]), .Cin(p_5_20[3]));
full_adder fa_6_20_1(.S(p_6_20[3]), .Cout(p_6_21[1]), .A(p_5_20[2]), .B(p_5_20[1]), .Cin(p_5_20[0]));
full_adder fa_6_21_0(.S(p_6_21[2]), .Cout(p_6_22[0]), .A(p_5_21[5]), .B(p_5_21[4]), .Cin(p_5_21[3]));
full_adder fa_6_21_1(.S(p_6_21[3]), .Cout(p_6_22[1]), .A(p_5_21[2]), .B(p_5_21[1]), .Cin(p_5_21[0]));
full_adder fa_6_22_0(.S(p_6_22[2]), .Cout(p_6_23[0]), .A(p_5_22[5]), .B(p_5_22[4]), .Cin(p_5_22[3]));
full_adder fa_6_22_1(.S(p_6_22[3]), .Cout(p_6_23[1]), .A(p_5_22[2]), .B(p_5_22[1]), .Cin(p_5_22[0]));
full_adder fa_6_23_0(.S(p_6_23[2]), .Cout(p_6_24[0]), .A(p_5_23[5]), .B(p_5_23[4]), .Cin(p_5_23[3]));
full_adder fa_6_23_1(.S(p_6_23[3]), .Cout(p_6_24[1]), .A(p_5_23[2]), .B(p_5_23[1]), .Cin(p_5_23[0]));
full_adder fa_6_24_0(.S(p_6_24[2]), .Cout(p_6_25[0]), .A(p_5_24[5]), .B(p_5_24[4]), .Cin(p_5_24[3]));
full_adder fa_6_24_1(.S(p_6_24[3]), .Cout(p_6_25[1]), .A(p_5_24[2]), .B(p_5_24[1]), .Cin(p_5_24[0]));
full_adder fa_6_25_0(.S(p_6_25[2]), .Cout(p_6_26[0]), .A(p_5_25[5]), .B(p_5_25[4]), .Cin(p_5_25[3]));
full_adder fa_6_25_1(.S(p_6_25[3]), .Cout(p_6_26[1]), .A(p_5_25[2]), .B(p_5_25[1]), .Cin(p_5_25[0]));
full_adder fa_6_26_0(.S(p_6_26[2]), .Cout(p_6_27[0]), .A(p_5_26[5]), .B(p_5_26[4]), .Cin(p_5_26[3]));
full_adder fa_6_26_1(.S(p_6_26[3]), .Cout(p_6_27[1]), .A(p_5_26[2]), .B(p_5_26[1]), .Cin(p_5_26[0]));
full_adder fa_6_27_0(.S(p_6_27[2]), .Cout(p_6_28[0]), .A(p_5_27[5]), .B(p_5_27[4]), .Cin(p_5_27[3]));
full_adder fa_6_27_1(.S(p_6_27[3]), .Cout(p_6_28[1]), .A(p_5_27[2]), .B(p_5_27[1]), .Cin(p_5_27[0]));
full_adder fa_6_28_0(.S(p_6_28[2]), .Cout(p_6_29[0]), .A(p_5_28[5]), .B(p_5_28[4]), .Cin(p_5_28[3]));
full_adder fa_6_28_1(.S(p_6_28[3]), .Cout(p_6_29[1]), .A(p_5_28[2]), .B(p_5_28[1]), .Cin(p_5_28[0]));
full_adder fa_6_29_0(.S(p_6_29[2]), .Cout(p_6_30[0]), .A(p_5_29[5]), .B(p_5_29[4]), .Cin(p_5_29[3]));
full_adder fa_6_29_1(.S(p_6_29[3]), .Cout(p_6_30[1]), .A(p_5_29[2]), .B(p_5_29[1]), .Cin(p_5_29[0]));
full_adder fa_6_30_0(.S(p_6_30[2]), .Cout(p_6_31[0]), .A(p_5_30[5]), .B(p_5_30[4]), .Cin(p_5_30[3]));
full_adder fa_6_30_1(.S(p_6_30[3]), .Cout(p_6_31[1]), .A(p_5_30[2]), .B(p_5_30[1]), .Cin(p_5_30[0]));
full_adder fa_6_31_0(.S(p_6_31[2]), .Cout(p_6_32[0]), .A(p_5_31[5]), .B(p_5_31[4]), .Cin(p_5_31[3]));
full_adder fa_6_31_1(.S(p_6_31[3]), .Cout(p_6_32[1]), .A(p_5_31[2]), .B(p_5_31[1]), .Cin(p_5_31[0]));
full_adder fa_6_32_0(.S(p_6_32[2]), .Cout(p_6_33[0]), .A(p_5_32[5]), .B(p_5_32[4]), .Cin(p_5_32[3]));
full_adder fa_6_32_1(.S(p_6_32[3]), .Cout(p_6_33[1]), .A(p_5_32[2]), .B(p_5_32[1]), .Cin(p_5_32[0]));
full_adder fa_6_33_0(.S(p_6_33[2]), .Cout(p_6_34[0]), .A(p_5_33[5]), .B(p_5_33[4]), .Cin(p_5_33[3]));
full_adder fa_6_33_1(.S(p_6_33[3]), .Cout(p_6_34[1]), .A(p_5_33[2]), .B(p_5_33[1]), .Cin(p_5_33[0]));
full_adder fa_6_34_0(.S(p_6_34[2]), .Cout(p_6_35[0]), .A(p_5_34[5]), .B(p_5_34[4]), .Cin(p_5_34[3]));
full_adder fa_6_34_1(.S(p_6_34[3]), .Cout(p_6_35[1]), .A(p_5_34[2]), .B(p_5_34[1]), .Cin(p_5_34[0]));
full_adder fa_6_35_0(.S(p_6_35[2]), .Cout(p_6_36[0]), .A(p_5_35[5]), .B(p_5_35[4]), .Cin(p_5_35[3]));
full_adder fa_6_35_1(.S(p_6_35[3]), .Cout(p_6_36[1]), .A(p_5_35[2]), .B(p_5_35[1]), .Cin(p_5_35[0]));
full_adder fa_6_36_0(.S(p_6_36[2]), .Cout(p_6_37[0]), .A(p_5_36[5]), .B(p_5_36[4]), .Cin(p_5_36[3]));
full_adder fa_6_36_1(.S(p_6_36[3]), .Cout(p_6_37[1]), .A(p_5_36[2]), .B(p_5_36[1]), .Cin(p_5_36[0]));
full_adder fa_6_37_0(.S(p_6_37[2]), .Cout(p_6_38[0]), .A(p_5_37[5]), .B(p_5_37[4]), .Cin(p_5_37[3]));
full_adder fa_6_37_1(.S(p_6_37[3]), .Cout(p_6_38[1]), .A(p_5_37[2]), .B(p_5_37[1]), .Cin(p_5_37[0]));
full_adder fa_6_38_0(.S(p_6_38[2]), .Cout(p_6_39[0]), .A(p_5_38[5]), .B(p_5_38[4]), .Cin(p_5_38[3]));
full_adder fa_6_38_1(.S(p_6_38[3]), .Cout(p_6_39[1]), .A(p_5_38[2]), .B(p_5_38[1]), .Cin(p_5_38[0]));
full_adder fa_6_39_0(.S(p_6_39[2]), .Cout(p_6_40[0]), .A(p_5_39[5]), .B(p_5_39[4]), .Cin(p_5_39[3]));
full_adder fa_6_39_1(.S(p_6_39[3]), .Cout(p_6_40[1]), .A(p_5_39[2]), .B(p_5_39[1]), .Cin(p_5_39[0]));
full_adder fa_6_40_0(.S(p_6_40[2]), .Cout(p_6_41[0]), .A(p_5_40[5]), .B(p_5_40[4]), .Cin(p_5_40[3]));
full_adder fa_6_40_1(.S(p_6_40[3]), .Cout(p_6_41[1]), .A(p_5_40[2]), .B(p_5_40[1]), .Cin(p_5_40[0]));
full_adder fa_6_41_0(.S(p_6_41[2]), .Cout(p_6_42[0]), .A(p_5_41[5]), .B(p_5_41[4]), .Cin(p_5_41[3]));
full_adder fa_6_41_1(.S(p_6_41[3]), .Cout(p_6_42[1]), .A(p_5_41[2]), .B(p_5_41[1]), .Cin(p_5_41[0]));
full_adder fa_6_42_0(.S(p_6_42[2]), .Cout(p_6_43[0]), .A(p_5_42[5]), .B(p_5_42[4]), .Cin(p_5_42[3]));
full_adder fa_6_42_1(.S(p_6_42[3]), .Cout(p_6_43[1]), .A(p_5_42[2]), .B(p_5_42[1]), .Cin(p_5_42[0]));
full_adder fa_6_43_0(.S(p_6_43[2]), .Cout(p_6_44[0]), .A(p_5_43[5]), .B(p_5_43[4]), .Cin(p_5_43[3]));
full_adder fa_6_43_1(.S(p_6_43[3]), .Cout(p_6_44[1]), .A(p_5_43[2]), .B(p_5_43[1]), .Cin(p_5_43[0]));
full_adder fa_6_44_0(.S(p_6_44[2]), .Cout(p_6_45[0]), .A(p_5_44[5]), .B(p_5_44[4]), .Cin(p_5_44[3]));
full_adder fa_6_44_1(.S(p_6_44[3]), .Cout(p_6_45[1]), .A(p_5_44[2]), .B(p_5_44[1]), .Cin(p_5_44[0]));
full_adder fa_6_45_0(.S(p_6_45[2]), .Cout(p_6_46[0]), .A(p_5_45[5]), .B(p_5_45[4]), .Cin(p_5_45[3]));
full_adder fa_6_45_1(.S(p_6_45[3]), .Cout(p_6_46[1]), .A(p_5_45[2]), .B(p_5_45[1]), .Cin(p_5_45[0]));
full_adder fa_6_46_0(.S(p_6_46[2]), .Cout(p_6_47[0]), .A(p_5_46[5]), .B(p_5_46[4]), .Cin(p_5_46[3]));
full_adder fa_6_46_1(.S(p_6_46[3]), .Cout(p_6_47[1]), .A(p_5_46[2]), .B(p_5_46[1]), .Cin(p_5_46[0]));
full_adder fa_6_47_0(.S(p_6_47[2]), .Cout(p_6_48[0]), .A(p_5_47[5]), .B(p_5_47[4]), .Cin(p_5_47[3]));
full_adder fa_6_47_1(.S(p_6_47[3]), .Cout(p_6_48[1]), .A(p_5_47[2]), .B(p_5_47[1]), .Cin(p_5_47[0]));
full_adder fa_6_48_0(.S(p_6_48[2]), .Cout(p_6_49[0]), .A(p_5_48[5]), .B(p_5_48[4]), .Cin(p_5_48[3]));
full_adder fa_6_48_1(.S(p_6_48[3]), .Cout(p_6_49[1]), .A(p_5_48[2]), .B(p_5_48[1]), .Cin(p_5_48[0]));
full_adder fa_6_49_0(.S(p_6_49[2]), .Cout(p_6_50[0]), .A(p_5_49[5]), .B(p_5_49[4]), .Cin(p_5_49[3]));
full_adder fa_6_49_1(.S(p_6_49[3]), .Cout(p_6_50[1]), .A(p_5_49[2]), .B(p_5_49[1]), .Cin(p_5_49[0]));
full_adder fa_6_50_0(.S(p_6_50[2]), .Cout(p_6_51[0]), .A(p_5_50[5]), .B(p_5_50[4]), .Cin(p_5_50[3]));
full_adder fa_6_50_1(.S(p_6_50[3]), .Cout(p_6_51[1]), .A(p_5_50[2]), .B(p_5_50[1]), .Cin(p_5_50[0]));
full_adder fa_6_51_0(.S(p_6_51[2]), .Cout(p_6_52[0]), .A(p_5_51[5]), .B(p_5_51[4]), .Cin(p_5_51[3]));
full_adder fa_6_51_1(.S(p_6_51[3]), .Cout(p_6_52[1]), .A(p_5_51[2]), .B(p_5_51[1]), .Cin(p_5_51[0]));
full_adder fa_6_52_0(.S(p_6_52[2]), .Cout(p_6_53[0]), .A(p_5_52[5]), .B(p_5_52[4]), .Cin(p_5_52[3]));
full_adder fa_6_52_1(.S(p_6_52[3]), .Cout(p_6_53[1]), .A(p_5_52[2]), .B(p_5_52[1]), .Cin(p_5_52[0]));
full_adder fa_6_53_0(.S(p_6_53[2]), .Cout(p_6_54[0]), .A(p_5_53[5]), .B(p_5_53[4]), .Cin(p_5_53[3]));
full_adder fa_6_53_1(.S(p_6_53[3]), .Cout(p_6_54[1]), .A(p_5_53[2]), .B(p_5_53[1]), .Cin(p_5_53[0]));
full_adder fa_6_54_0(.S(p_6_54[2]), .Cout(p_6_55[0]), .A(p_5_54[5]), .B(p_5_54[4]), .Cin(p_5_54[3]));
full_adder fa_6_54_1(.S(p_6_54[3]), .Cout(p_6_55[1]), .A(p_5_54[2]), .B(p_5_54[1]), .Cin(p_5_54[0]));
full_adder fa_6_55_0(.S(p_6_55[2]), .Cout(p_6_56[0]), .A(p_5_55[5]), .B(p_5_55[4]), .Cin(p_5_55[3]));
full_adder fa_6_55_1(.S(p_6_55[3]), .Cout(p_6_56[1]), .A(p_5_55[2]), .B(p_5_55[1]), .Cin(p_5_55[0]));
full_adder fa_6_56_0(.S(p_6_56[2]), .Cout(p_6_57[0]), .A(p_5_56[5]), .B(p_5_56[4]), .Cin(p_5_56[3]));
full_adder fa_6_56_1(.S(p_6_56[3]), .Cout(p_6_57[1]), .A(p_5_56[2]), .B(p_5_56[1]), .Cin(p_5_56[0]));
full_adder fa_6_57_0(.S(p_6_57[2]), .Cout(p_6_58[0]), .A(p_5_57[5]), .B(p_5_57[4]), .Cin(p_5_57[3]));
full_adder fa_6_57_1(.S(p_6_57[3]), .Cout(p_6_58[1]), .A(p_5_57[2]), .B(p_5_57[1]), .Cin(p_5_57[0]));
full_adder fa_6_58_0(.S(p_6_58[2]), .Cout(p_6_59[0]), .A(p_5_58[5]), .B(p_5_58[4]), .Cin(p_5_58[3]));
full_adder fa_6_58_1(.S(p_6_58[3]), .Cout(p_6_59[1]), .A(p_5_58[2]), .B(p_5_58[1]), .Cin(p_5_58[0]));
full_adder fa_6_59_0(.S(p_6_59[2]), .Cout(p_6_60[0]), .A(p_5_59[3]), .B(p_5_59[2]), .Cin(p_5_59[1]));

// Stage 7 non-added partial products
assign p_7_0[0:0] = p_6_0[0:0];
assign p_7_1[1:0] = p_6_1[1:0];
assign p_7_2[2:0] = p_6_2[2:0];
assign p_7_3[2:1] = p_6_3[1:0];
assign p_7_4[2:2] = p_6_4[0:0];
assign p_7_5[2:2] = p_6_5[0:0];
assign p_7_6[2:2] = p_6_6[0:0];
assign p_7_7[2:2] = p_6_7[0:0];
assign p_7_8[2:2] = p_6_8[0:0];
assign p_7_9[2:2] = p_6_9[0:0];
assign p_7_10[2:2] = p_6_10[0:0];
assign p_7_11[2:2] = p_6_11[0:0];
assign p_7_12[2:2] = p_6_12[0:0];
assign p_7_13[2:2] = p_6_13[0:0];
assign p_7_14[2:2] = p_6_14[0:0];
assign p_7_15[2:2] = p_6_15[0:0];
assign p_7_16[2:2] = p_6_16[0:0];
assign p_7_17[2:2] = p_6_17[0:0];
assign p_7_18[2:2] = p_6_18[0:0];
assign p_7_19[2:2] = p_6_19[0:0];
assign p_7_20[2:2] = p_6_20[0:0];
assign p_7_21[2:2] = p_6_21[0:0];
assign p_7_22[2:2] = p_6_22[0:0];
assign p_7_23[2:2] = p_6_23[0:0];
assign p_7_24[2:2] = p_6_24[0:0];
assign p_7_25[2:2] = p_6_25[0:0];
assign p_7_26[2:2] = p_6_26[0:0];
assign p_7_27[2:2] = p_6_27[0:0];
assign p_7_28[2:2] = p_6_28[0:0];
assign p_7_29[2:2] = p_6_29[0:0];
assign p_7_30[2:2] = p_6_30[0:0];
assign p_7_31[2:2] = p_6_31[0:0];
assign p_7_32[2:2] = p_6_32[0:0];
assign p_7_33[2:2] = p_6_33[0:0];
assign p_7_34[2:2] = p_6_34[0:0];
assign p_7_35[2:2] = p_6_35[0:0];
assign p_7_36[2:2] = p_6_36[0:0];
assign p_7_37[2:2] = p_6_37[0:0];
assign p_7_38[2:2] = p_6_38[0:0];
assign p_7_39[2:2] = p_6_39[0:0];
assign p_7_40[2:2] = p_6_40[0:0];
assign p_7_41[2:2] = p_6_41[0:0];
assign p_7_42[2:2] = p_6_42[0:0];
assign p_7_43[2:2] = p_6_43[0:0];
assign p_7_44[2:2] = p_6_44[0:0];
assign p_7_45[2:2] = p_6_45[0:0];
assign p_7_46[2:2] = p_6_46[0:0];
assign p_7_47[2:2] = p_6_47[0:0];
assign p_7_48[2:2] = p_6_48[0:0];
assign p_7_49[2:2] = p_6_49[0:0];
assign p_7_50[2:2] = p_6_50[0:0];
assign p_7_51[2:2] = p_6_51[0:0];
assign p_7_52[2:2] = p_6_52[0:0];
assign p_7_53[2:2] = p_6_53[0:0];
assign p_7_54[2:2] = p_6_54[0:0];
assign p_7_55[2:2] = p_6_55[0:0];
assign p_7_56[2:2] = p_6_56[0:0];
assign p_7_57[2:2] = p_6_57[0:0];
assign p_7_58[2:2] = p_6_58[0:0];
assign p_7_59[2:2] = p_6_59[0:0];
assign p_7_60[2:2] = p_6_60[0:0];
assign p_7_61[2:1] = p_6_61[1:0];
assign p_7_62[0:0] = p_6_62[0:0];
// Stage 7 adders
half_adder ha_7_3(.S(p_7_3[0]), .Cout(p_7_4[0]), .A(p_6_3[3]), .B(p_6_3[2]));
full_adder fa_7_4_0(.S(p_7_4[1]), .Cout(p_7_5[0]), .A(p_6_4[3]), .B(p_6_4[2]), .Cin(p_6_4[1]));
full_adder fa_7_5_0(.S(p_7_5[1]), .Cout(p_7_6[0]), .A(p_6_5[3]), .B(p_6_5[2]), .Cin(p_6_5[1]));
full_adder fa_7_6_0(.S(p_7_6[1]), .Cout(p_7_7[0]), .A(p_6_6[3]), .B(p_6_6[2]), .Cin(p_6_6[1]));
full_adder fa_7_7_0(.S(p_7_7[1]), .Cout(p_7_8[0]), .A(p_6_7[3]), .B(p_6_7[2]), .Cin(p_6_7[1]));
full_adder fa_7_8_0(.S(p_7_8[1]), .Cout(p_7_9[0]), .A(p_6_8[3]), .B(p_6_8[2]), .Cin(p_6_8[1]));
full_adder fa_7_9_0(.S(p_7_9[1]), .Cout(p_7_10[0]), .A(p_6_9[3]), .B(p_6_9[2]), .Cin(p_6_9[1]));
full_adder fa_7_10_0(.S(p_7_10[1]), .Cout(p_7_11[0]), .A(p_6_10[3]), .B(p_6_10[2]), .Cin(p_6_10[1]));
full_adder fa_7_11_0(.S(p_7_11[1]), .Cout(p_7_12[0]), .A(p_6_11[3]), .B(p_6_11[2]), .Cin(p_6_11[1]));
full_adder fa_7_12_0(.S(p_7_12[1]), .Cout(p_7_13[0]), .A(p_6_12[3]), .B(p_6_12[2]), .Cin(p_6_12[1]));
full_adder fa_7_13_0(.S(p_7_13[1]), .Cout(p_7_14[0]), .A(p_6_13[3]), .B(p_6_13[2]), .Cin(p_6_13[1]));
full_adder fa_7_14_0(.S(p_7_14[1]), .Cout(p_7_15[0]), .A(p_6_14[3]), .B(p_6_14[2]), .Cin(p_6_14[1]));
full_adder fa_7_15_0(.S(p_7_15[1]), .Cout(p_7_16[0]), .A(p_6_15[3]), .B(p_6_15[2]), .Cin(p_6_15[1]));
full_adder fa_7_16_0(.S(p_7_16[1]), .Cout(p_7_17[0]), .A(p_6_16[3]), .B(p_6_16[2]), .Cin(p_6_16[1]));
full_adder fa_7_17_0(.S(p_7_17[1]), .Cout(p_7_18[0]), .A(p_6_17[3]), .B(p_6_17[2]), .Cin(p_6_17[1]));
full_adder fa_7_18_0(.S(p_7_18[1]), .Cout(p_7_19[0]), .A(p_6_18[3]), .B(p_6_18[2]), .Cin(p_6_18[1]));
full_adder fa_7_19_0(.S(p_7_19[1]), .Cout(p_7_20[0]), .A(p_6_19[3]), .B(p_6_19[2]), .Cin(p_6_19[1]));
full_adder fa_7_20_0(.S(p_7_20[1]), .Cout(p_7_21[0]), .A(p_6_20[3]), .B(p_6_20[2]), .Cin(p_6_20[1]));
full_adder fa_7_21_0(.S(p_7_21[1]), .Cout(p_7_22[0]), .A(p_6_21[3]), .B(p_6_21[2]), .Cin(p_6_21[1]));
full_adder fa_7_22_0(.S(p_7_22[1]), .Cout(p_7_23[0]), .A(p_6_22[3]), .B(p_6_22[2]), .Cin(p_6_22[1]));
full_adder fa_7_23_0(.S(p_7_23[1]), .Cout(p_7_24[0]), .A(p_6_23[3]), .B(p_6_23[2]), .Cin(p_6_23[1]));
full_adder fa_7_24_0(.S(p_7_24[1]), .Cout(p_7_25[0]), .A(p_6_24[3]), .B(p_6_24[2]), .Cin(p_6_24[1]));
full_adder fa_7_25_0(.S(p_7_25[1]), .Cout(p_7_26[0]), .A(p_6_25[3]), .B(p_6_25[2]), .Cin(p_6_25[1]));
full_adder fa_7_26_0(.S(p_7_26[1]), .Cout(p_7_27[0]), .A(p_6_26[3]), .B(p_6_26[2]), .Cin(p_6_26[1]));
full_adder fa_7_27_0(.S(p_7_27[1]), .Cout(p_7_28[0]), .A(p_6_27[3]), .B(p_6_27[2]), .Cin(p_6_27[1]));
full_adder fa_7_28_0(.S(p_7_28[1]), .Cout(p_7_29[0]), .A(p_6_28[3]), .B(p_6_28[2]), .Cin(p_6_28[1]));
full_adder fa_7_29_0(.S(p_7_29[1]), .Cout(p_7_30[0]), .A(p_6_29[3]), .B(p_6_29[2]), .Cin(p_6_29[1]));
full_adder fa_7_30_0(.S(p_7_30[1]), .Cout(p_7_31[0]), .A(p_6_30[3]), .B(p_6_30[2]), .Cin(p_6_30[1]));
full_adder fa_7_31_0(.S(p_7_31[1]), .Cout(p_7_32[0]), .A(p_6_31[3]), .B(p_6_31[2]), .Cin(p_6_31[1]));
full_adder fa_7_32_0(.S(p_7_32[1]), .Cout(p_7_33[0]), .A(p_6_32[3]), .B(p_6_32[2]), .Cin(p_6_32[1]));
full_adder fa_7_33_0(.S(p_7_33[1]), .Cout(p_7_34[0]), .A(p_6_33[3]), .B(p_6_33[2]), .Cin(p_6_33[1]));
full_adder fa_7_34_0(.S(p_7_34[1]), .Cout(p_7_35[0]), .A(p_6_34[3]), .B(p_6_34[2]), .Cin(p_6_34[1]));
full_adder fa_7_35_0(.S(p_7_35[1]), .Cout(p_7_36[0]), .A(p_6_35[3]), .B(p_6_35[2]), .Cin(p_6_35[1]));
full_adder fa_7_36_0(.S(p_7_36[1]), .Cout(p_7_37[0]), .A(p_6_36[3]), .B(p_6_36[2]), .Cin(p_6_36[1]));
full_adder fa_7_37_0(.S(p_7_37[1]), .Cout(p_7_38[0]), .A(p_6_37[3]), .B(p_6_37[2]), .Cin(p_6_37[1]));
full_adder fa_7_38_0(.S(p_7_38[1]), .Cout(p_7_39[0]), .A(p_6_38[3]), .B(p_6_38[2]), .Cin(p_6_38[1]));
full_adder fa_7_39_0(.S(p_7_39[1]), .Cout(p_7_40[0]), .A(p_6_39[3]), .B(p_6_39[2]), .Cin(p_6_39[1]));
full_adder fa_7_40_0(.S(p_7_40[1]), .Cout(p_7_41[0]), .A(p_6_40[3]), .B(p_6_40[2]), .Cin(p_6_40[1]));
full_adder fa_7_41_0(.S(p_7_41[1]), .Cout(p_7_42[0]), .A(p_6_41[3]), .B(p_6_41[2]), .Cin(p_6_41[1]));
full_adder fa_7_42_0(.S(p_7_42[1]), .Cout(p_7_43[0]), .A(p_6_42[3]), .B(p_6_42[2]), .Cin(p_6_42[1]));
full_adder fa_7_43_0(.S(p_7_43[1]), .Cout(p_7_44[0]), .A(p_6_43[3]), .B(p_6_43[2]), .Cin(p_6_43[1]));
full_adder fa_7_44_0(.S(p_7_44[1]), .Cout(p_7_45[0]), .A(p_6_44[3]), .B(p_6_44[2]), .Cin(p_6_44[1]));
full_adder fa_7_45_0(.S(p_7_45[1]), .Cout(p_7_46[0]), .A(p_6_45[3]), .B(p_6_45[2]), .Cin(p_6_45[1]));
full_adder fa_7_46_0(.S(p_7_46[1]), .Cout(p_7_47[0]), .A(p_6_46[3]), .B(p_6_46[2]), .Cin(p_6_46[1]));
full_adder fa_7_47_0(.S(p_7_47[1]), .Cout(p_7_48[0]), .A(p_6_47[3]), .B(p_6_47[2]), .Cin(p_6_47[1]));
full_adder fa_7_48_0(.S(p_7_48[1]), .Cout(p_7_49[0]), .A(p_6_48[3]), .B(p_6_48[2]), .Cin(p_6_48[1]));
full_adder fa_7_49_0(.S(p_7_49[1]), .Cout(p_7_50[0]), .A(p_6_49[3]), .B(p_6_49[2]), .Cin(p_6_49[1]));
full_adder fa_7_50_0(.S(p_7_50[1]), .Cout(p_7_51[0]), .A(p_6_50[3]), .B(p_6_50[2]), .Cin(p_6_50[1]));
full_adder fa_7_51_0(.S(p_7_51[1]), .Cout(p_7_52[0]), .A(p_6_51[3]), .B(p_6_51[2]), .Cin(p_6_51[1]));
full_adder fa_7_52_0(.S(p_7_52[1]), .Cout(p_7_53[0]), .A(p_6_52[3]), .B(p_6_52[2]), .Cin(p_6_52[1]));
full_adder fa_7_53_0(.S(p_7_53[1]), .Cout(p_7_54[0]), .A(p_6_53[3]), .B(p_6_53[2]), .Cin(p_6_53[1]));
full_adder fa_7_54_0(.S(p_7_54[1]), .Cout(p_7_55[0]), .A(p_6_54[3]), .B(p_6_54[2]), .Cin(p_6_54[1]));
full_adder fa_7_55_0(.S(p_7_55[1]), .Cout(p_7_56[0]), .A(p_6_55[3]), .B(p_6_55[2]), .Cin(p_6_55[1]));
full_adder fa_7_56_0(.S(p_7_56[1]), .Cout(p_7_57[0]), .A(p_6_56[3]), .B(p_6_56[2]), .Cin(p_6_56[1]));
full_adder fa_7_57_0(.S(p_7_57[1]), .Cout(p_7_58[0]), .A(p_6_57[3]), .B(p_6_57[2]), .Cin(p_6_57[1]));
full_adder fa_7_58_0(.S(p_7_58[1]), .Cout(p_7_59[0]), .A(p_6_58[3]), .B(p_6_58[2]), .Cin(p_6_58[1]));
full_adder fa_7_59_0(.S(p_7_59[1]), .Cout(p_7_60[0]), .A(p_6_59[3]), .B(p_6_59[2]), .Cin(p_6_59[1]));
full_adder fa_7_60_0(.S(p_7_60[1]), .Cout(p_7_61[0]), .A(p_6_60[3]), .B(p_6_60[2]), .Cin(p_6_60[1]));

// Stage 8 non-added partial products
assign p_8_0[0:0] = p_7_0[0:0];
assign p_8_1[1:0] = p_7_1[1:0];
assign p_8_2[1:1] = p_7_2[0:0];
assign p_8_62[1:1] = p_7_62[0:0];
// Stage 8 adders
half_adder ha_8_2(.S(p_8_2[0]), .Cout(p_8_3[0]), .A(p_7_2[2]), .B(p_7_2[1]));
full_adder fa_8_3_0(.S(p_8_3[1]), .Cout(p_8_4[0]), .A(p_7_3[2]), .B(p_7_3[1]), .Cin(p_7_3[0]));
full_adder fa_8_4_0(.S(p_8_4[1]), .Cout(p_8_5[0]), .A(p_7_4[2]), .B(p_7_4[1]), .Cin(p_7_4[0]));
full_adder fa_8_5_0(.S(p_8_5[1]), .Cout(p_8_6[0]), .A(p_7_5[2]), .B(p_7_5[1]), .Cin(p_7_5[0]));
full_adder fa_8_6_0(.S(p_8_6[1]), .Cout(p_8_7[0]), .A(p_7_6[2]), .B(p_7_6[1]), .Cin(p_7_6[0]));
full_adder fa_8_7_0(.S(p_8_7[1]), .Cout(p_8_8[0]), .A(p_7_7[2]), .B(p_7_7[1]), .Cin(p_7_7[0]));
full_adder fa_8_8_0(.S(p_8_8[1]), .Cout(p_8_9[0]), .A(p_7_8[2]), .B(p_7_8[1]), .Cin(p_7_8[0]));
full_adder fa_8_9_0(.S(p_8_9[1]), .Cout(p_8_10[0]), .A(p_7_9[2]), .B(p_7_9[1]), .Cin(p_7_9[0]));
full_adder fa_8_10_0(.S(p_8_10[1]), .Cout(p_8_11[0]), .A(p_7_10[2]), .B(p_7_10[1]), .Cin(p_7_10[0]));
full_adder fa_8_11_0(.S(p_8_11[1]), .Cout(p_8_12[0]), .A(p_7_11[2]), .B(p_7_11[1]), .Cin(p_7_11[0]));
full_adder fa_8_12_0(.S(p_8_12[1]), .Cout(p_8_13[0]), .A(p_7_12[2]), .B(p_7_12[1]), .Cin(p_7_12[0]));
full_adder fa_8_13_0(.S(p_8_13[1]), .Cout(p_8_14[0]), .A(p_7_13[2]), .B(p_7_13[1]), .Cin(p_7_13[0]));
full_adder fa_8_14_0(.S(p_8_14[1]), .Cout(p_8_15[0]), .A(p_7_14[2]), .B(p_7_14[1]), .Cin(p_7_14[0]));
full_adder fa_8_15_0(.S(p_8_15[1]), .Cout(p_8_16[0]), .A(p_7_15[2]), .B(p_7_15[1]), .Cin(p_7_15[0]));
full_adder fa_8_16_0(.S(p_8_16[1]), .Cout(p_8_17[0]), .A(p_7_16[2]), .B(p_7_16[1]), .Cin(p_7_16[0]));
full_adder fa_8_17_0(.S(p_8_17[1]), .Cout(p_8_18[0]), .A(p_7_17[2]), .B(p_7_17[1]), .Cin(p_7_17[0]));
full_adder fa_8_18_0(.S(p_8_18[1]), .Cout(p_8_19[0]), .A(p_7_18[2]), .B(p_7_18[1]), .Cin(p_7_18[0]));
full_adder fa_8_19_0(.S(p_8_19[1]), .Cout(p_8_20[0]), .A(p_7_19[2]), .B(p_7_19[1]), .Cin(p_7_19[0]));
full_adder fa_8_20_0(.S(p_8_20[1]), .Cout(p_8_21[0]), .A(p_7_20[2]), .B(p_7_20[1]), .Cin(p_7_20[0]));
full_adder fa_8_21_0(.S(p_8_21[1]), .Cout(p_8_22[0]), .A(p_7_21[2]), .B(p_7_21[1]), .Cin(p_7_21[0]));
full_adder fa_8_22_0(.S(p_8_22[1]), .Cout(p_8_23[0]), .A(p_7_22[2]), .B(p_7_22[1]), .Cin(p_7_22[0]));
full_adder fa_8_23_0(.S(p_8_23[1]), .Cout(p_8_24[0]), .A(p_7_23[2]), .B(p_7_23[1]), .Cin(p_7_23[0]));
full_adder fa_8_24_0(.S(p_8_24[1]), .Cout(p_8_25[0]), .A(p_7_24[2]), .B(p_7_24[1]), .Cin(p_7_24[0]));
full_adder fa_8_25_0(.S(p_8_25[1]), .Cout(p_8_26[0]), .A(p_7_25[2]), .B(p_7_25[1]), .Cin(p_7_25[0]));
full_adder fa_8_26_0(.S(p_8_26[1]), .Cout(p_8_27[0]), .A(p_7_26[2]), .B(p_7_26[1]), .Cin(p_7_26[0]));
full_adder fa_8_27_0(.S(p_8_27[1]), .Cout(p_8_28[0]), .A(p_7_27[2]), .B(p_7_27[1]), .Cin(p_7_27[0]));
full_adder fa_8_28_0(.S(p_8_28[1]), .Cout(p_8_29[0]), .A(p_7_28[2]), .B(p_7_28[1]), .Cin(p_7_28[0]));
full_adder fa_8_29_0(.S(p_8_29[1]), .Cout(p_8_30[0]), .A(p_7_29[2]), .B(p_7_29[1]), .Cin(p_7_29[0]));
full_adder fa_8_30_0(.S(p_8_30[1]), .Cout(p_8_31[0]), .A(p_7_30[2]), .B(p_7_30[1]), .Cin(p_7_30[0]));
full_adder fa_8_31_0(.S(p_8_31[1]), .Cout(p_8_32[0]), .A(p_7_31[2]), .B(p_7_31[1]), .Cin(p_7_31[0]));
full_adder fa_8_32_0(.S(p_8_32[1]), .Cout(p_8_33[0]), .A(p_7_32[2]), .B(p_7_32[1]), .Cin(p_7_32[0]));
full_adder fa_8_33_0(.S(p_8_33[1]), .Cout(p_8_34[0]), .A(p_7_33[2]), .B(p_7_33[1]), .Cin(p_7_33[0]));
full_adder fa_8_34_0(.S(p_8_34[1]), .Cout(p_8_35[0]), .A(p_7_34[2]), .B(p_7_34[1]), .Cin(p_7_34[0]));
full_adder fa_8_35_0(.S(p_8_35[1]), .Cout(p_8_36[0]), .A(p_7_35[2]), .B(p_7_35[1]), .Cin(p_7_35[0]));
full_adder fa_8_36_0(.S(p_8_36[1]), .Cout(p_8_37[0]), .A(p_7_36[2]), .B(p_7_36[1]), .Cin(p_7_36[0]));
full_adder fa_8_37_0(.S(p_8_37[1]), .Cout(p_8_38[0]), .A(p_7_37[2]), .B(p_7_37[1]), .Cin(p_7_37[0]));
full_adder fa_8_38_0(.S(p_8_38[1]), .Cout(p_8_39[0]), .A(p_7_38[2]), .B(p_7_38[1]), .Cin(p_7_38[0]));
full_adder fa_8_39_0(.S(p_8_39[1]), .Cout(p_8_40[0]), .A(p_7_39[2]), .B(p_7_39[1]), .Cin(p_7_39[0]));
full_adder fa_8_40_0(.S(p_8_40[1]), .Cout(p_8_41[0]), .A(p_7_40[2]), .B(p_7_40[1]), .Cin(p_7_40[0]));
full_adder fa_8_41_0(.S(p_8_41[1]), .Cout(p_8_42[0]), .A(p_7_41[2]), .B(p_7_41[1]), .Cin(p_7_41[0]));
full_adder fa_8_42_0(.S(p_8_42[1]), .Cout(p_8_43[0]), .A(p_7_42[2]), .B(p_7_42[1]), .Cin(p_7_42[0]));
full_adder fa_8_43_0(.S(p_8_43[1]), .Cout(p_8_44[0]), .A(p_7_43[2]), .B(p_7_43[1]), .Cin(p_7_43[0]));
full_adder fa_8_44_0(.S(p_8_44[1]), .Cout(p_8_45[0]), .A(p_7_44[2]), .B(p_7_44[1]), .Cin(p_7_44[0]));
full_adder fa_8_45_0(.S(p_8_45[1]), .Cout(p_8_46[0]), .A(p_7_45[2]), .B(p_7_45[1]), .Cin(p_7_45[0]));
full_adder fa_8_46_0(.S(p_8_46[1]), .Cout(p_8_47[0]), .A(p_7_46[2]), .B(p_7_46[1]), .Cin(p_7_46[0]));
full_adder fa_8_47_0(.S(p_8_47[1]), .Cout(p_8_48[0]), .A(p_7_47[2]), .B(p_7_47[1]), .Cin(p_7_47[0]));
full_adder fa_8_48_0(.S(p_8_48[1]), .Cout(p_8_49[0]), .A(p_7_48[2]), .B(p_7_48[1]), .Cin(p_7_48[0]));
full_adder fa_8_49_0(.S(p_8_49[1]), .Cout(p_8_50[0]), .A(p_7_49[2]), .B(p_7_49[1]), .Cin(p_7_49[0]));
full_adder fa_8_50_0(.S(p_8_50[1]), .Cout(p_8_51[0]), .A(p_7_50[2]), .B(p_7_50[1]), .Cin(p_7_50[0]));
full_adder fa_8_51_0(.S(p_8_51[1]), .Cout(p_8_52[0]), .A(p_7_51[2]), .B(p_7_51[1]), .Cin(p_7_51[0]));
full_adder fa_8_52_0(.S(p_8_52[1]), .Cout(p_8_53[0]), .A(p_7_52[2]), .B(p_7_52[1]), .Cin(p_7_52[0]));
full_adder fa_8_53_0(.S(p_8_53[1]), .Cout(p_8_54[0]), .A(p_7_53[2]), .B(p_7_53[1]), .Cin(p_7_53[0]));
full_adder fa_8_54_0(.S(p_8_54[1]), .Cout(p_8_55[0]), .A(p_7_54[2]), .B(p_7_54[1]), .Cin(p_7_54[0]));
full_adder fa_8_55_0(.S(p_8_55[1]), .Cout(p_8_56[0]), .A(p_7_55[2]), .B(p_7_55[1]), .Cin(p_7_55[0]));
full_adder fa_8_56_0(.S(p_8_56[1]), .Cout(p_8_57[0]), .A(p_7_56[2]), .B(p_7_56[1]), .Cin(p_7_56[0]));
full_adder fa_8_57_0(.S(p_8_57[1]), .Cout(p_8_58[0]), .A(p_7_57[2]), .B(p_7_57[1]), .Cin(p_7_57[0]));
full_adder fa_8_58_0(.S(p_8_58[1]), .Cout(p_8_59[0]), .A(p_7_58[2]), .B(p_7_58[1]), .Cin(p_7_58[0]));
full_adder fa_8_59_0(.S(p_8_59[1]), .Cout(p_8_60[0]), .A(p_7_59[2]), .B(p_7_59[1]), .Cin(p_7_59[0]));
full_adder fa_8_60_0(.S(p_8_60[1]), .Cout(p_8_61[0]), .A(p_7_60[2]), .B(p_7_60[1]), .Cin(p_7_60[0]));
full_adder fa_8_61_0(.S(p_8_61[1]), .Cout(p_8_62[0]), .A(p_7_61[2]), .B(p_7_61[1]), .Cin(p_7_61[0]));

// Final stage
wire [63:0] f1;
wire [63:0] f2;
assign f1 = {1'b0, p_8_61[0], p_8_60[0], p_8_59[0], p_8_58[0], p_8_57[0], p_8_56[0], p_8_55[0], p_8_54[0], p_8_53[0], p_8_52[0], p_8_51[0], p_8_50[0], p_8_49[0], p_8_48[0], p_8_47[0], p_8_46[0], p_8_45[0], p_8_44[0], p_8_43[0], p_8_42[0], p_8_41[0], p_8_40[0], p_8_39[0], p_8_38[0], p_8_37[0], p_8_36[0], p_8_35[0], p_8_34[0], p_8_33[0], p_8_32[0], p_8_31[0], p_8_30[0], p_8_29[0], p_8_28[0], p_8_27[0], p_8_26[0], p_8_25[0], p_8_24[0], p_8_23[0], p_8_22[0], p_8_21[0], p_8_20[0], p_8_19[0], p_8_18[0], p_8_17[0], p_8_16[0], p_8_15[0], p_8_14[0], p_8_13[0], p_8_12[0], p_8_11[0], p_8_10[0], p_8_9[0], p_8_8[0], p_8_7[0], p_8_6[0], p_8_5[0], p_8_4[0], p_8_3[0], p_8_2[0], p_8_1[0], p_8_0[0]};
assign f2 = {1'b0, p_8_61[1], p_8_60[1], p_8_59[1], p_8_58[1], p_8_57[1], p_8_56[1], p_8_55[1], p_8_54[1], p_8_53[1], p_8_52[1], p_8_51[1], p_8_50[1], p_8_49[1], p_8_48[1], p_8_47[1], p_8_46[1], p_8_45[1], p_8_44[1], p_8_43[1], p_8_42[1], p_8_41[1], p_8_40[1], p_8_39[1], p_8_38[1], p_8_37[1], p_8_36[1], p_8_35[1], p_8_34[1], p_8_33[1], p_8_32[1], p_8_31[1], p_8_30[1], p_8_29[1], p_8_28[1], p_8_27[1], p_8_26[1], p_8_25[1], p_8_24[1], p_8_23[1], p_8_22[1], p_8_21[1], p_8_20[1], p_8_19[1], p_8_18[1], p_8_17[1], p_8_16[1], p_8_15[1], p_8_14[1], p_8_13[1], p_8_12[1], p_8_11[1], p_8_10[1], p_8_9[1], p_8_8[1], p_8_7[1], p_8_6[1], p_8_5[1], p_8_4[1], p_8_3[1], p_8_2[1], p_8_1[1], 1'b0};
// Insert final adder
cla_64 cla(.A(f1), .B(f2), .Cin(1'b0), .Sum(Product));
endmodule
