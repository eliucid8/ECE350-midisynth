module midibuffer(
    output[7:0] msg, input sig, input clock);
    
endmodule